
module bootrom(addr_i_2_, addr_i_3_, addr_i_4_, addr_i_5_, addr_i_6_, addr_i_7_, addr_i_8_, addr_i_9_, addr_i_10_, addr_i_11_, addr_i_12_, data_o_0_, data_o_1_
, data_o_2_, data_o_3_, data_o_4_, data_o_5_, data_o_6_, data_o_7_, data_o_8_, data_o_9_, data_o_10_, data_o_11_, data_o_12_, data_o_13_, data_o_14_, data_o_15_, data_o_16_, data_o_17_, data_o_18_, data_o_19_, data_o_20_, data_o_21_, data_o_22_
, data_o_23_, data_o_24_, data_o_25_, data_o_26_, data_o_27_, data_o_28_, data_o_29_, data_o_30_, data_o_31_);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  input addr_i_10_;
  wire addr_i_10_;
  input addr_i_11_;
  wire addr_i_11_;
  input addr_i_12_;
  wire addr_i_12_;
  input addr_i_2_;
  wire addr_i_2_;
  input addr_i_3_;
  wire addr_i_3_;
  input addr_i_4_;
  wire addr_i_4_;
  input addr_i_5_;
  wire addr_i_5_;
  input addr_i_6_;
  wire addr_i_6_;
  input addr_i_7_;
  wire addr_i_7_;
  input addr_i_8_;
  wire addr_i_8_;
  input addr_i_9_;
  wire addr_i_9_;
  output data_o_0_;
  wire data_o_0_;
  output data_o_10_;
  wire data_o_10_;
  output data_o_11_;
  wire data_o_11_;
  output data_o_12_;
  wire data_o_12_;
  output data_o_13_;
  wire data_o_13_;
  output data_o_14_;
  wire data_o_14_;
  output data_o_15_;
  wire data_o_15_;
  output data_o_16_;
  wire data_o_16_;
  output data_o_17_;
  wire data_o_17_;
  output data_o_18_;
  wire data_o_18_;
  output data_o_19_;
  wire data_o_19_;
  output data_o_1_;
  wire data_o_1_;
  output data_o_20_;
  wire data_o_20_;
  output data_o_21_;
  wire data_o_21_;
  output data_o_22_;
  wire data_o_22_;
  output data_o_23_;
  wire data_o_23_;
  output data_o_24_;
  wire data_o_24_;
  output data_o_25_;
  wire data_o_25_;
  output data_o_26_;
  wire data_o_26_;
  output data_o_27_;
  wire data_o_27_;
  output data_o_28_;
  wire data_o_28_;
  output data_o_29_;
  wire data_o_29_;
  output data_o_2_;
  wire data_o_2_;
  output data_o_30_;
  wire data_o_30_;
  output data_o_31_;
  wire data_o_31_;
  output data_o_3_;
  wire data_o_3_;
  output data_o_4_;
  wire data_o_4_;
  output data_o_5_;
  wire data_o_5_;
  output data_o_6_;
  wire data_o_6_;
  output data_o_7_;
  wire data_o_7_;
  output data_o_8_;
  wire data_o_8_;
  output data_o_9_;
  wire data_o_9_;
  sg13g2_inv_1 _09514_ (
    .A(addr_i_10_),
    .Y(_03731_)
  );
  sg13g2_buf_1 _09515_ (
    .A(_03731_),
    .X(_03841_)
  );
  sg13g2_nand2_1 _09516_ (
    .A(addr_i_4_),
    .B(addr_i_5_),
    .Y(_03952_)
  );
  sg13g2_buf_1 _09517_ (
    .A(_03952_),
    .X(_04063_)
  );
  sg13g2_nor2b_1 _09518_ (
    .A(addr_i_6_),
    .B_N(addr_i_7_),
    .Y(_04173_)
  );
  sg13g2_buf_1 _09519_ (
    .A(_04173_),
    .X(_04284_)
  );
  sg13g2_or3_1 _09520_ (
    .A(addr_i_4_),
    .B(addr_i_7_),
    .C(addr_i_5_),
    .X(_04395_)
  );
  sg13g2_o21ai_1 _09521_ (
    .A1(_04063_),
    .A2(_04284_),
    .B1(_04395_),
    .Y(_04505_)
  );
  sg13g2_nand2_1 _09522_ (
    .A(addr_i_6_),
    .B(addr_i_5_),
    .Y(_04616_)
  );
  sg13g2_or2_1 _09523_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .X(_04726_)
  );
  sg13g2_nor2_1 _09524_ (
    .A(_04616_),
    .B(_04726_),
    .Y(_04837_)
  );
  sg13g2_a21o_1 _09525_ (
    .A1(addr_i_2_),
    .A2(_04505_),
    .B1(_04837_),
    .X(_04948_)
  );
  sg13g2_and2_1 _09526_ (
    .A(addr_i_7_),
    .B(addr_i_5_),
    .X(_05058_)
  );
  sg13g2_buf_1 _09527_ (
    .A(_05058_),
    .X(_05169_)
  );
  sg13g2_buf_1 _09528_ (
    .A(_05169_),
    .X(_05280_)
  );
  sg13g2_nor2b_1 _09529_ (
    .A(addr_i_4_),
    .B_N(addr_i_2_),
    .Y(_05390_)
  );
  sg13g2_buf_1 _09530_ (
    .A(_05390_),
    .X(_05501_)
  );
  sg13g2_nand2_1 _09531_ (
    .A(_05280_),
    .B(_05501_),
    .Y(_05611_)
  );
  sg13g2_nor2_1 _09532_ (
    .A(addr_i_7_),
    .B(addr_i_5_),
    .Y(_05722_)
  );
  sg13g2_buf_1 _09533_ (
    .A(_05722_),
    .X(_05833_)
  );
  sg13g2_nor2_1 _09534_ (
    .A(addr_i_3_),
    .B(addr_i_2_),
    .Y(_05943_)
  );
  sg13g2_buf_1 _09535_ (
    .A(_05943_),
    .X(_06054_)
  );
  sg13g2_nand2_1 _09536_ (
    .A(_05833_),
    .B(_06054_),
    .Y(_06164_)
  );
  sg13g2_inv_1 _09537_ (
    .A(addr_i_6_),
    .Y(_06275_)
  );
  sg13g2_buf_1 _09538_ (
    .A(_06275_),
    .X(_06386_)
  );
  sg13g2_buf_1 _09539_ (
    .A(_06386_),
    .X(_06496_)
  );
  sg13g2_buf_1 _09540_ (
    .A(_06496_),
    .X(_06607_)
  );
  sg13g2_buf_1 _09541_ (
    .A(_06607_),
    .X(_06717_)
  );
  sg13g2_a21oi_1 _09542_ (
    .A1(_05611_),
    .A2(_06164_),
    .B1(_06717_),
    .Y(_06828_)
  );
  sg13g2_inv_1 _09543_ (
    .A(addr_i_3_),
    .Y(_06938_)
  );
  sg13g2_buf_1 _09544_ (
    .A(_06938_),
    .X(_07049_)
  );
  sg13g2_nor2b_1 _09545_ (
    .A(addr_i_2_),
    .B_N(addr_i_5_),
    .Y(_07159_)
  );
  sg13g2_nor2_1 _09546_ (
    .A(_07049_),
    .B(_07159_),
    .Y(_07270_)
  );
  sg13g2_inv_1 _09547_ (
    .A(addr_i_2_),
    .Y(_07381_)
  );
  sg13g2_buf_1 _09548_ (
    .A(_07381_),
    .X(_07491_)
  );
  sg13g2_nand2b_1 _09549_ (
    .A_N(addr_i_5_),
    .B(addr_i_7_),
    .Y(_07602_)
  );
  sg13g2_nor2_1 _09550_ (
    .A(_07491_),
    .B(_07602_),
    .Y(_07712_)
  );
  sg13g2_inv_1 _09551_ (
    .A(addr_i_4_),
    .Y(_07823_)
  );
  sg13g2_buf_1 _09552_ (
    .A(_07823_),
    .X(_07933_)
  );
  sg13g2_buf_1 _09553_ (
    .A(_07933_),
    .X(_08044_)
  );
  sg13g2_buf_1 _09554_ (
    .A(_08044_),
    .X(_08155_)
  );
  sg13g2_o21ai_1 _09555_ (
    .A1(_07270_),
    .A2(_07712_),
    .B1(_08155_),
    .Y(_08265_)
  );
  sg13g2_buf_1 _09556_ (
    .A(_07602_),
    .X(_08376_)
  );
  sg13g2_nand2_1 _09557_ (
    .A(addr_i_4_),
    .B(_08376_),
    .Y(_08486_)
  );
  sg13g2_nor2b_1 _09558_ (
    .A(addr_i_5_),
    .B_N(addr_i_7_),
    .Y(_08597_)
  );
  sg13g2_nand2_1 _09559_ (
    .A(addr_i_3_),
    .B(_08597_),
    .Y(_08707_)
  );
  sg13g2_o21ai_1 _09560_ (
    .A1(addr_i_3_),
    .A2(_08486_),
    .B1(_08707_),
    .Y(_08818_)
  );
  sg13g2_nand2b_1 _09561_ (
    .A_N(addr_i_7_),
    .B(addr_i_4_),
    .Y(_08929_)
  );
  sg13g2_buf_1 _09562_ (
    .A(_06938_),
    .X(_09038_)
  );
  sg13g2_nand2_1 _09563_ (
    .A(_09038_),
    .B(_05169_),
    .Y(_09149_)
  );
  sg13g2_a21oi_1 _09564_ (
    .A1(_08929_),
    .A2(_09149_),
    .B1(addr_i_2_),
    .Y(_09259_)
  );
  sg13g2_nor2_1 _09565_ (
    .A(_08818_),
    .B(_09259_),
    .Y(_09370_)
  );
  sg13g2_a21oi_1 _09566_ (
    .A1(_08265_),
    .A2(_09370_),
    .B1(addr_i_6_),
    .Y(_09470_)
  );
  sg13g2_a22oi_1 _09567_ (
    .A1(addr_i_3_),
    .A2(_04948_),
    .B1(_06828_),
    .B2(_09470_),
    .Y(_09481_)
  );
  sg13g2_buf_1 _09568_ (
    .A(_08929_),
    .X(_09492_)
  );
  sg13g2_and2_1 _09569_ (
    .A(addr_i_6_),
    .B(addr_i_5_),
    .X(_09503_)
  );
  sg13g2_buf_1 _09570_ (
    .A(_09503_),
    .X(_00000_)
  );
  sg13g2_buf_1 _09571_ (
    .A(_00000_),
    .X(_00011_)
  );
  sg13g2_buf_1 _09572_ (
    .A(_00011_),
    .X(_00022_)
  );
  sg13g2_buf_1 _09573_ (
    .A(_07823_),
    .X(_00033_)
  );
  sg13g2_buf_1 _09574_ (
    .A(_00033_),
    .X(_00044_)
  );
  sg13g2_nand2_1 _09575_ (
    .A(_00044_),
    .B(_05169_),
    .Y(_00055_)
  );
  sg13g2_nor2b_1 _09576_ (
    .A(addr_i_7_),
    .B_N(addr_i_6_),
    .Y(_00066_)
  );
  sg13g2_nand2_1 _09577_ (
    .A(addr_i_4_),
    .B(_00066_),
    .Y(_00077_)
  );
  sg13g2_a21o_1 _09578_ (
    .A1(_00055_),
    .A2(_00077_),
    .B1(addr_i_3_),
    .X(_00088_)
  );
  sg13g2_nor2_1 _09579_ (
    .A(addr_i_4_),
    .B(addr_i_7_),
    .Y(_00099_)
  );
  sg13g2_buf_1 _09580_ (
    .A(_00099_),
    .X(_00110_)
  );
  sg13g2_and3_1 _09581_ (
    .A(addr_i_4_),
    .B(addr_i_7_),
    .C(addr_i_6_),
    .X(_00121_)
  );
  sg13g2_buf_1 _09582_ (
    .A(_00121_),
    .X(_00132_)
  );
  sg13g2_o21ai_1 _09583_ (
    .A1(_00110_),
    .A2(_00132_),
    .B1(addr_i_3_),
    .Y(_00143_)
  );
  sg13g2_nor2b_1 _09584_ (
    .A(addr_i_7_),
    .B_N(addr_i_5_),
    .Y(_00154_)
  );
  sg13g2_buf_1 _09585_ (
    .A(_00154_),
    .X(_00165_)
  );
  sg13g2_inv_1 _09586_ (
    .A(addr_i_7_),
    .Y(_00176_)
  );
  sg13g2_or2_1 _09587_ (
    .A(addr_i_6_),
    .B(addr_i_5_),
    .X(_00187_)
  );
  sg13g2_buf_1 _09588_ (
    .A(_00187_),
    .X(_00198_)
  );
  sg13g2_nor2_1 _09589_ (
    .A(_00176_),
    .B(_00198_),
    .Y(_00209_)
  );
  sg13g2_o21ai_1 _09590_ (
    .A1(_00165_),
    .A2(_00209_),
    .B1(addr_i_4_),
    .Y(_00220_)
  );
  sg13g2_nor2_1 _09591_ (
    .A(addr_i_6_),
    .B(addr_i_5_),
    .Y(_00231_)
  );
  sg13g2_buf_1 _09592_ (
    .A(_00231_),
    .X(_00242_)
  );
  sg13g2_nand2_1 _09593_ (
    .A(_00110_),
    .B(_00242_),
    .Y(_00253_)
  );
  sg13g2_nand4_1 _09594_ (
    .A(_00088_),
    .B(_00143_),
    .C(_00220_),
    .D(_00253_),
    .Y(_00264_)
  );
  sg13g2_nor2_1 _09595_ (
    .A(addr_i_6_),
    .B(_05169_),
    .Y(_00275_)
  );
  sg13g2_nand2_1 _09596_ (
    .A(addr_i_3_),
    .B(_00275_),
    .Y(_00286_)
  );
  sg13g2_buf_1 _09597_ (
    .A(_08597_),
    .X(_00297_)
  );
  sg13g2_nor2_1 _09598_ (
    .A(addr_i_3_),
    .B(addr_i_4_),
    .Y(_00308_)
  );
  sg13g2_buf_1 _09599_ (
    .A(_00308_),
    .X(_00319_)
  );
  sg13g2_o21ai_1 _09600_ (
    .A1(addr_i_6_),
    .A2(_00297_),
    .B1(_00319_),
    .Y(_00330_)
  );
  sg13g2_a21oi_1 _09601_ (
    .A1(_00286_),
    .A2(_00330_),
    .B1(addr_i_2_),
    .Y(_00341_)
  );
  sg13g2_a221oi_1 _09602_ (
    .A1(_09492_),
    .A2(_00022_),
    .B1(_00264_),
    .B2(addr_i_2_),
    .C1(_00341_),
    .Y(_00352_)
  );
  sg13g2_nor2_1 _09603_ (
    .A(addr_i_8_),
    .B(_00352_),
    .Y(_00363_)
  );
  sg13g2_inv_1 _09604_ (
    .A(addr_i_9_),
    .Y(_00374_)
  );
  sg13g2_buf_1 _09605_ (
    .A(_00374_),
    .X(_00385_)
  );
  sg13g2_buf_1 _09606_ (
    .A(_00385_),
    .X(_00396_)
  );
  sg13g2_a22oi_1 _09607_ (
    .A1(addr_i_8_),
    .A2(_09481_),
    .B1(_00363_),
    .B2(_00396_),
    .Y(_00407_)
  );
  sg13g2_nor2_1 _09608_ (
    .A(addr_i_8_),
    .B(addr_i_7_),
    .Y(_00418_)
  );
  sg13g2_buf_1 _09609_ (
    .A(_00418_),
    .X(_00429_)
  );
  sg13g2_buf_1 _09610_ (
    .A(_00429_),
    .X(_00440_)
  );
  sg13g2_nand2b_1 _09611_ (
    .A_N(addr_i_2_),
    .B(addr_i_5_),
    .Y(_00451_)
  );
  sg13g2_buf_1 _09612_ (
    .A(_00451_),
    .X(_00462_)
  );
  sg13g2_nand2_1 _09613_ (
    .A(_06386_),
    .B(_00462_),
    .Y(_00473_)
  );
  sg13g2_buf_1 _09614_ (
    .A(_06386_),
    .X(_00484_)
  );
  sg13g2_xnor2_1 _09615_ (
    .A(addr_i_2_),
    .B(addr_i_5_),
    .Y(_00495_)
  );
  sg13g2_nand2_1 _09616_ (
    .A(_00484_),
    .B(_00495_),
    .Y(_00506_)
  );
  sg13g2_nor2_1 _09617_ (
    .A(addr_i_3_),
    .B(_00506_),
    .Y(_00517_)
  );
  sg13g2_a22oi_1 _09618_ (
    .A1(addr_i_3_),
    .A2(_00473_),
    .B1(_00517_),
    .B2(addr_i_4_),
    .Y(_00528_)
  );
  sg13g2_nor2b_1 _09619_ (
    .A(addr_i_6_),
    .B_N(addr_i_5_),
    .Y(_00539_)
  );
  sg13g2_buf_1 _09620_ (
    .A(_00539_),
    .X(_00550_)
  );
  sg13g2_buf_1 _09621_ (
    .A(_00550_),
    .X(_00561_)
  );
  sg13g2_and2_1 _09622_ (
    .A(addr_i_3_),
    .B(addr_i_2_),
    .X(_00572_)
  );
  sg13g2_buf_1 _09623_ (
    .A(_00572_),
    .X(_00583_)
  );
  sg13g2_buf_1 _09624_ (
    .A(_00583_),
    .X(_00594_)
  );
  sg13g2_nor2b_1 _09625_ (
    .A(addr_i_3_),
    .B_N(addr_i_6_),
    .Y(_00605_)
  );
  sg13g2_buf_1 _09626_ (
    .A(_00605_),
    .X(_00616_)
  );
  sg13g2_buf_1 _09627_ (
    .A(_00616_),
    .X(_00626_)
  );
  sg13g2_buf_1 _09628_ (
    .A(_00033_),
    .X(_00637_)
  );
  sg13g2_buf_1 _09629_ (
    .A(_00637_),
    .X(_00648_)
  );
  sg13g2_buf_1 _09630_ (
    .A(_00648_),
    .X(_00659_)
  );
  sg13g2_a22oi_1 _09631_ (
    .A1(_00561_),
    .A2(_00594_),
    .B1(_00626_),
    .B2(_00659_),
    .Y(_00670_)
  );
  sg13g2_or2_1 _09632_ (
    .A(addr_i_3_),
    .B(addr_i_2_),
    .X(_00681_)
  );
  sg13g2_buf_1 _09633_ (
    .A(_00681_),
    .X(_00692_)
  );
  sg13g2_buf_1 _09634_ (
    .A(_00692_),
    .X(_00703_)
  );
  sg13g2_nand2_1 _09635_ (
    .A(addr_i_2_),
    .B(addr_i_5_),
    .Y(_00714_)
  );
  sg13g2_buf_1 _09636_ (
    .A(_00714_),
    .X(_00725_)
  );
  sg13g2_buf_1 _09637_ (
    .A(_00725_),
    .X(_00736_)
  );
  sg13g2_buf_1 _09638_ (
    .A(_00736_),
    .X(_00747_)
  );
  sg13g2_nand3_1 _09639_ (
    .A(addr_i_6_),
    .B(_00703_),
    .C(_00747_),
    .Y(_00758_)
  );
  sg13g2_o21ai_1 _09640_ (
    .A1(_00528_),
    .A2(_00670_),
    .B1(_00758_),
    .Y(_00769_)
  );
  sg13g2_nand2b_1 _09641_ (
    .A_N(addr_i_8_),
    .B(addr_i_7_),
    .Y(_00780_)
  );
  sg13g2_buf_1 _09642_ (
    .A(_00780_),
    .X(_00791_)
  );
  sg13g2_buf_1 _09643_ (
    .A(_00791_),
    .X(_00802_)
  );
  sg13g2_nand2b_1 _09644_ (
    .A_N(addr_i_2_),
    .B(addr_i_3_),
    .Y(_00813_)
  );
  sg13g2_nor2_1 _09645_ (
    .A(_04616_),
    .B(_00813_),
    .Y(_00824_)
  );
  sg13g2_xor2_1 _09646_ (
    .A(addr_i_6_),
    .B(addr_i_5_),
    .X(_00835_)
  );
  sg13g2_nand2_1 _09647_ (
    .A(addr_i_2_),
    .B(_00835_),
    .Y(_00846_)
  );
  sg13g2_nor2_1 _09648_ (
    .A(addr_i_3_),
    .B(_00846_),
    .Y(_00857_)
  );
  sg13g2_nor3_1 _09649_ (
    .A(addr_i_4_),
    .B(_00824_),
    .C(_00857_),
    .Y(_00868_)
  );
  sg13g2_nor2_1 _09650_ (
    .A(addr_i_2_),
    .B(addr_i_6_),
    .Y(_00879_)
  );
  sg13g2_buf_1 _09651_ (
    .A(_00879_),
    .X(_00890_)
  );
  sg13g2_nor2_1 _09652_ (
    .A(addr_i_5_),
    .B(_00890_),
    .Y(_00901_)
  );
  sg13g2_nand2b_1 _09653_ (
    .A_N(addr_i_6_),
    .B(addr_i_5_),
    .Y(_00912_)
  );
  sg13g2_buf_1 _09654_ (
    .A(_00912_),
    .X(_00923_)
  );
  sg13g2_nor2_1 _09655_ (
    .A(addr_i_2_),
    .B(_00923_),
    .Y(_00934_)
  );
  sg13g2_buf_1 _09656_ (
    .A(_00934_),
    .X(_00945_)
  );
  sg13g2_buf_1 _09657_ (
    .A(_00044_),
    .X(_00956_)
  );
  sg13g2_buf_1 _09658_ (
    .A(_00956_),
    .X(_00967_)
  );
  sg13g2_a22oi_1 _09659_ (
    .A1(addr_i_3_),
    .A2(_00901_),
    .B1(_00945_),
    .B2(_00967_),
    .Y(_00978_)
  );
  sg13g2_nor2_1 _09660_ (
    .A(_00868_),
    .B(_00978_),
    .Y(_00989_)
  );
  sg13g2_nand2_1 _09661_ (
    .A(addr_i_8_),
    .B(addr_i_7_),
    .Y(_01000_)
  );
  sg13g2_buf_1 _09662_ (
    .A(_01000_),
    .X(_01011_)
  );
  sg13g2_nor2b_1 _09663_ (
    .A(addr_i_4_),
    .B_N(addr_i_6_),
    .Y(_01022_)
  );
  sg13g2_buf_1 _09664_ (
    .A(_01022_),
    .X(_01033_)
  );
  sg13g2_nor2_1 _09665_ (
    .A(addr_i_5_),
    .B(_01033_),
    .Y(_01044_)
  );
  sg13g2_nand2b_1 _09666_ (
    .A_N(addr_i_6_),
    .B(addr_i_2_),
    .Y(_01055_)
  );
  sg13g2_buf_1 _09667_ (
    .A(_01055_),
    .X(_01066_)
  );
  sg13g2_buf_1 _09668_ (
    .A(_01066_),
    .X(_01077_)
  );
  sg13g2_nand2_1 _09669_ (
    .A(_00033_),
    .B(_07159_),
    .Y(_01087_)
  );
  sg13g2_a21oi_1 _09670_ (
    .A1(_01077_),
    .A2(_01087_),
    .B1(addr_i_3_),
    .Y(_01098_)
  );
  sg13g2_nor4_1 _09671_ (
    .A(_01011_),
    .B(_01044_),
    .C(_00824_),
    .D(_01098_),
    .Y(_01109_)
  );
  sg13g2_buf_1 _09672_ (
    .A(_00044_),
    .X(_01120_)
  );
  sg13g2_buf_1 _09673_ (
    .A(_01120_),
    .X(_01131_)
  );
  sg13g2_and2_1 _09674_ (
    .A(addr_i_2_),
    .B(addr_i_5_),
    .X(_01142_)
  );
  sg13g2_buf_1 _09675_ (
    .A(_01142_),
    .X(_01153_)
  );
  sg13g2_nor2_1 _09676_ (
    .A(_01153_),
    .B(_00890_),
    .Y(_01164_)
  );
  sg13g2_nand2_1 _09677_ (
    .A(_07491_),
    .B(_00539_),
    .Y(_01175_)
  );
  sg13g2_o21ai_1 _09678_ (
    .A1(addr_i_3_),
    .A2(_01164_),
    .B1(_01175_),
    .Y(_01186_)
  );
  sg13g2_nand2b_1 _09679_ (
    .A_N(addr_i_5_),
    .B(addr_i_3_),
    .Y(_01197_)
  );
  sg13g2_buf_1 _09680_ (
    .A(_01197_),
    .X(_01208_)
  );
  sg13g2_nand2_1 _09681_ (
    .A(_07049_),
    .B(_07159_),
    .Y(_01219_)
  );
  sg13g2_buf_1 _09682_ (
    .A(_01219_),
    .X(_01230_)
  );
  sg13g2_nand2_1 _09683_ (
    .A(addr_i_4_),
    .B(addr_i_6_),
    .Y(_01241_)
  );
  sg13g2_buf_1 _09684_ (
    .A(_01241_),
    .X(_01252_)
  );
  sg13g2_a21oi_1 _09685_ (
    .A1(_01208_),
    .A2(_01230_),
    .B1(_01252_),
    .Y(_01263_)
  );
  sg13g2_nand2_1 _09686_ (
    .A(addr_i_8_),
    .B(_00176_),
    .Y(_01274_)
  );
  sg13g2_buf_1 _09687_ (
    .A(_01274_),
    .X(_01285_)
  );
  sg13g2_a22oi_1 _09688_ (
    .A1(_01131_),
    .A2(_01186_),
    .B1(_01263_),
    .B2(_01285_),
    .Y(_01296_)
  );
  sg13g2_nor3_1 _09689_ (
    .A(addr_i_9_),
    .B(_01109_),
    .C(_01296_),
    .Y(_01307_)
  );
  sg13g2_o21ai_1 _09690_ (
    .A1(_00802_),
    .A2(_00989_),
    .B1(_01307_),
    .Y(_01318_)
  );
  sg13g2_a21oi_1 _09691_ (
    .A1(_00440_),
    .A2(_00769_),
    .B1(_01318_),
    .Y(_01329_)
  );
  sg13g2_nor3_1 _09692_ (
    .A(_03841_),
    .B(_00407_),
    .C(_01329_),
    .Y(_01340_)
  );
  sg13g2_buf_1 _09693_ (
    .A(_00385_),
    .X(_01351_)
  );
  sg13g2_or2_1 _09694_ (
    .A(addr_i_2_),
    .B(addr_i_5_),
    .X(_01362_)
  );
  sg13g2_buf_1 _09695_ (
    .A(_01362_),
    .X(_01373_)
  );
  sg13g2_buf_1 _09696_ (
    .A(_01373_),
    .X(_01384_)
  );
  sg13g2_nand3b_1 _09697_ (
    .A_N(addr_i_6_),
    .B(addr_i_5_),
    .C(addr_i_2_),
    .Y(_01395_)
  );
  sg13g2_buf_1 _09698_ (
    .A(_01395_),
    .X(_01406_)
  );
  sg13g2_a21oi_1 _09699_ (
    .A1(_01384_),
    .A2(_01406_),
    .B1(addr_i_3_),
    .Y(_01417_)
  );
  sg13g2_o21ai_1 _09700_ (
    .A1(_00824_),
    .A2(_01417_),
    .B1(addr_i_4_),
    .Y(_01428_)
  );
  sg13g2_and2_1 _09701_ (
    .A(addr_i_3_),
    .B(addr_i_6_),
    .X(_01439_)
  );
  sg13g2_buf_1 _09702_ (
    .A(_01439_),
    .X(_01450_)
  );
  sg13g2_nor2b_1 _09703_ (
    .A(addr_i_2_),
    .B_N(addr_i_4_),
    .Y(_01461_)
  );
  sg13g2_buf_1 _09704_ (
    .A(_01461_),
    .X(_01472_)
  );
  sg13g2_nor2_1 _09705_ (
    .A(addr_i_5_),
    .B(_01472_),
    .Y(_01483_)
  );
  sg13g2_buf_1 _09706_ (
    .A(_01274_),
    .X(_01494_)
  );
  sg13g2_a21oi_1 _09707_ (
    .A1(_01450_),
    .A2(_01483_),
    .B1(_01494_),
    .Y(_01505_)
  );
  sg13g2_nand2_1 _09708_ (
    .A(_01428_),
    .B(_01505_),
    .Y(_01515_)
  );
  sg13g2_inv_1 _09709_ (
    .A(addr_i_8_),
    .Y(_01526_)
  );
  sg13g2_buf_1 _09710_ (
    .A(_01526_),
    .X(_01537_)
  );
  sg13g2_buf_1 _09711_ (
    .A(_01537_),
    .X(_01548_)
  );
  sg13g2_buf_1 _09712_ (
    .A(_01548_),
    .X(_01559_)
  );
  sg13g2_buf_1 _09713_ (
    .A(_00198_),
    .X(_01570_)
  );
  sg13g2_buf_1 _09714_ (
    .A(_04616_),
    .X(_01581_)
  );
  sg13g2_or2_1 _09715_ (
    .A(addr_i_2_),
    .B(addr_i_7_),
    .X(_01592_)
  );
  sg13g2_buf_1 _09716_ (
    .A(_01592_),
    .X(_01603_)
  );
  sg13g2_a22oi_1 _09717_ (
    .A1(_01570_),
    .A2(_01581_),
    .B1(addr_i_4_),
    .B2(_01603_),
    .Y(_01614_)
  );
  sg13g2_nand2b_1 _09718_ (
    .A_N(addr_i_5_),
    .B(addr_i_4_),
    .Y(_01625_)
  );
  sg13g2_buf_1 _09719_ (
    .A(_01625_),
    .X(_01636_)
  );
  sg13g2_nand3b_1 _09720_ (
    .A_N(addr_i_7_),
    .B(addr_i_6_),
    .C(addr_i_2_),
    .Y(_01647_)
  );
  sg13g2_buf_1 _09721_ (
    .A(_01647_),
    .X(_01658_)
  );
  sg13g2_and2_1 _09722_ (
    .A(addr_i_7_),
    .B(addr_i_6_),
    .X(_01669_)
  );
  sg13g2_buf_1 _09723_ (
    .A(_01669_),
    .X(_01680_)
  );
  sg13g2_nand2_1 _09724_ (
    .A(_01680_),
    .B(_05390_),
    .Y(_01691_)
  );
  sg13g2_o21ai_1 _09725_ (
    .A1(_01636_),
    .A2(_01658_),
    .B1(_01691_),
    .Y(_01702_)
  );
  sg13g2_o21ai_1 _09726_ (
    .A1(_01614_),
    .A2(_01702_),
    .B1(addr_i_3_),
    .Y(_01713_)
  );
  sg13g2_or2_1 _09727_ (
    .A(addr_i_3_),
    .B(addr_i_4_),
    .X(_01724_)
  );
  sg13g2_nor2_1 _09728_ (
    .A(_00451_),
    .B(_01724_),
    .Y(_01735_)
  );
  sg13g2_buf_1 _09729_ (
    .A(_01735_),
    .X(_01746_)
  );
  sg13g2_buf_1 _09730_ (
    .A(_00198_),
    .X(_01757_)
  );
  sg13g2_nand3b_1 _09731_ (
    .A_N(addr_i_2_),
    .B(addr_i_6_),
    .C(addr_i_5_),
    .Y(_01768_)
  );
  sg13g2_a21oi_1 _09732_ (
    .A1(_01757_),
    .A2(_01768_),
    .B1(_08044_),
    .Y(_01779_)
  );
  sg13g2_o21ai_1 _09733_ (
    .A1(_01746_),
    .A2(_01779_),
    .B1(addr_i_7_),
    .Y(_01790_)
  );
  sg13g2_nand3_1 _09734_ (
    .A(_01559_),
    .B(_01713_),
    .C(_01790_),
    .Y(_01801_)
  );
  sg13g2_nand2_1 _09735_ (
    .A(_01515_),
    .B(_01801_),
    .Y(_01812_)
  );
  sg13g2_nand3b_1 _09736_ (
    .A_N(addr_i_5_),
    .B(addr_i_2_),
    .C(addr_i_4_),
    .Y(_01823_)
  );
  sg13g2_buf_1 _09737_ (
    .A(_01823_),
    .X(_01834_)
  );
  sg13g2_a21oi_1 _09738_ (
    .A1(_01834_),
    .A2(_01087_),
    .B1(addr_i_3_),
    .Y(_01845_)
  );
  sg13g2_nor2_1 _09739_ (
    .A(addr_i_7_),
    .B(addr_i_6_),
    .Y(_01856_)
  );
  sg13g2_buf_1 _09740_ (
    .A(_01856_),
    .X(_01867_)
  );
  sg13g2_buf_1 _09741_ (
    .A(_01867_),
    .X(_01878_)
  );
  sg13g2_buf_1 _09742_ (
    .A(_05390_),
    .X(_01888_)
  );
  sg13g2_nand2b_1 _09743_ (
    .A_N(addr_i_2_),
    .B(addr_i_4_),
    .Y(_01899_)
  );
  sg13g2_nor2_1 _09744_ (
    .A(addr_i_5_),
    .B(_01899_),
    .Y(_01910_)
  );
  sg13g2_o21ai_1 _09745_ (
    .A1(_01888_),
    .A2(_01910_),
    .B1(addr_i_3_),
    .Y(_01921_)
  );
  sg13g2_nand3b_1 _09746_ (
    .A_N(_01845_),
    .B(_01878_),
    .C(_01921_),
    .Y(_01932_)
  );
  sg13g2_and2_1 _09747_ (
    .A(addr_i_3_),
    .B(addr_i_5_),
    .X(_01943_)
  );
  sg13g2_buf_1 _09748_ (
    .A(_01943_),
    .X(_01954_)
  );
  sg13g2_nand2_1 _09749_ (
    .A(addr_i_2_),
    .B(addr_i_6_),
    .Y(_01965_)
  );
  sg13g2_buf_1 _09750_ (
    .A(_01965_),
    .X(_01976_)
  );
  sg13g2_nand2_1 _09751_ (
    .A(_00033_),
    .B(_00879_),
    .Y(_01987_)
  );
  sg13g2_nand2_1 _09752_ (
    .A(_01976_),
    .B(_01987_),
    .Y(_01998_)
  );
  sg13g2_nand2b_1 _09753_ (
    .A_N(addr_i_5_),
    .B(addr_i_6_),
    .Y(_02009_)
  );
  sg13g2_buf_1 _09754_ (
    .A(_02009_),
    .X(_02020_)
  );
  sg13g2_buf_1 _09755_ (
    .A(_04726_),
    .X(_02031_)
  );
  sg13g2_nor2_1 _09756_ (
    .A(_02020_),
    .B(_02031_),
    .Y(_02042_)
  );
  sg13g2_buf_1 _09757_ (
    .A(_00176_),
    .X(_02053_)
  );
  sg13g2_buf_1 _09758_ (
    .A(_02053_),
    .X(_02064_)
  );
  sg13g2_a22oi_1 _09759_ (
    .A1(_01954_),
    .A2(_01998_),
    .B1(_02042_),
    .B2(_02064_),
    .Y(_02075_)
  );
  sg13g2_buf_1 _09760_ (
    .A(_07049_),
    .X(_02086_)
  );
  sg13g2_nor2b_1 _09761_ (
    .A(addr_i_5_),
    .B_N(addr_i_6_),
    .Y(_02097_)
  );
  sg13g2_buf_1 _09762_ (
    .A(_02097_),
    .X(_02108_)
  );
  sg13g2_nor2_1 _09763_ (
    .A(addr_i_2_),
    .B(_02108_),
    .Y(_02119_)
  );
  sg13g2_nor2_1 _09764_ (
    .A(_02086_),
    .B(_02119_),
    .Y(_02130_)
  );
  sg13g2_buf_1 _09765_ (
    .A(_01142_),
    .X(_02141_)
  );
  sg13g2_buf_1 _09766_ (
    .A(_02097_),
    .X(_02152_)
  );
  sg13g2_nor3_1 _09767_ (
    .A(addr_i_3_),
    .B(_02141_),
    .C(_02152_),
    .Y(_02163_)
  );
  sg13g2_o21ai_1 _09768_ (
    .A1(_02130_),
    .A2(_02163_),
    .B1(addr_i_4_),
    .Y(_02174_)
  );
  sg13g2_nand2b_1 _09769_ (
    .A_N(addr_i_3_),
    .B(addr_i_2_),
    .Y(_02185_)
  );
  sg13g2_buf_1 _09770_ (
    .A(_02185_),
    .X(_02196_)
  );
  sg13g2_nand2_1 _09771_ (
    .A(addr_i_3_),
    .B(addr_i_5_),
    .Y(_02207_)
  );
  sg13g2_buf_1 _09772_ (
    .A(_02207_),
    .X(_02218_)
  );
  sg13g2_nand2_1 _09773_ (
    .A(_02196_),
    .B(_02218_),
    .Y(_02229_)
  );
  sg13g2_or3_1 _09774_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .C(addr_i_5_),
    .X(_02240_)
  );
  sg13g2_buf_1 _09775_ (
    .A(_02240_),
    .X(_02250_)
  );
  sg13g2_a21oi_1 _09776_ (
    .A1(_00725_),
    .A2(_02250_),
    .B1(addr_i_3_),
    .Y(_02261_)
  );
  sg13g2_nand2b_1 _09777_ (
    .A_N(addr_i_7_),
    .B(addr_i_6_),
    .Y(_02272_)
  );
  sg13g2_buf_1 _09778_ (
    .A(_02272_),
    .X(_02283_)
  );
  sg13g2_buf_1 _09779_ (
    .A(_02283_),
    .X(_02294_)
  );
  sg13g2_a22oi_1 _09780_ (
    .A1(addr_i_4_),
    .A2(_02229_),
    .B1(_02261_),
    .B2(_02294_),
    .Y(_02305_)
  );
  sg13g2_a22oi_1 _09781_ (
    .A1(_02075_),
    .A2(_02174_),
    .B1(_02305_),
    .B2(addr_i_8_),
    .Y(_02316_)
  );
  sg13g2_nor2_1 _09782_ (
    .A(_08044_),
    .B(_08376_),
    .Y(_02327_)
  );
  sg13g2_nand3b_1 _09783_ (
    .A_N(addr_i_2_),
    .B(addr_i_7_),
    .C(addr_i_5_),
    .Y(_02338_)
  );
  sg13g2_buf_1 _09784_ (
    .A(_02338_),
    .X(_02349_)
  );
  sg13g2_nand2_1 _09785_ (
    .A(addr_i_7_),
    .B(addr_i_5_),
    .Y(_02360_)
  );
  sg13g2_buf_1 _09786_ (
    .A(_02360_),
    .X(_02371_)
  );
  sg13g2_nand2_1 _09787_ (
    .A(addr_i_2_),
    .B(_02371_),
    .Y(_02382_)
  );
  sg13g2_a21oi_1 _09788_ (
    .A1(_02349_),
    .A2(_02382_),
    .B1(addr_i_4_),
    .Y(_02393_)
  );
  sg13g2_buf_1 _09789_ (
    .A(_02086_),
    .X(_02404_)
  );
  sg13g2_o21ai_1 _09790_ (
    .A1(_02327_),
    .A2(_02393_),
    .B1(_02404_),
    .Y(_02415_)
  );
  sg13g2_xnor2_1 _09791_ (
    .A(addr_i_7_),
    .B(addr_i_6_),
    .Y(_02426_)
  );
  sg13g2_buf_1 _09792_ (
    .A(_02426_),
    .X(_02437_)
  );
  sg13g2_a21oi_1 _09793_ (
    .A1(_00637_),
    .A2(_08597_),
    .B1(_00154_),
    .Y(_02448_)
  );
  sg13g2_buf_1 _09794_ (
    .A(_00813_),
    .X(_02459_)
  );
  sg13g2_buf_1 _09795_ (
    .A(_02459_),
    .X(_02470_)
  );
  sg13g2_a21oi_1 _09796_ (
    .A1(_08486_),
    .A2(_02448_),
    .B1(_02470_),
    .Y(_02481_)
  );
  sg13g2_nor2_1 _09797_ (
    .A(_02437_),
    .B(_02481_),
    .Y(_02492_)
  );
  sg13g2_nor2b_1 _09798_ (
    .A(addr_i_5_),
    .B_N(addr_i_3_),
    .Y(_02503_)
  );
  sg13g2_buf_1 _09799_ (
    .A(_02503_),
    .X(_02514_)
  );
  sg13g2_xnor2_1 _09800_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .Y(_02525_)
  );
  sg13g2_buf_1 _09801_ (
    .A(_02525_),
    .X(_02536_)
  );
  sg13g2_or2_1 _09802_ (
    .A(addr_i_7_),
    .B(addr_i_6_),
    .X(_02547_)
  );
  sg13g2_buf_1 _09803_ (
    .A(_02547_),
    .X(_02558_)
  );
  sg13g2_buf_1 _09804_ (
    .A(_02558_),
    .X(_02569_)
  );
  sg13g2_a22oi_1 _09805_ (
    .A1(_02514_),
    .A2(_02536_),
    .B1(_01746_),
    .B2(_02569_),
    .Y(_02580_)
  );
  sg13g2_nand2b_1 _09806_ (
    .A_N(addr_i_4_),
    .B(addr_i_5_),
    .Y(_02591_)
  );
  sg13g2_buf_1 _09807_ (
    .A(_02591_),
    .X(_02602_)
  );
  sg13g2_a21oi_1 _09808_ (
    .A1(addr_i_2_),
    .A2(_02602_),
    .B1(addr_i_3_),
    .Y(_02613_)
  );
  sg13g2_buf_1 _09809_ (
    .A(_01669_),
    .X(_02623_)
  );
  sg13g2_buf_1 _09810_ (
    .A(_01625_),
    .X(_02634_)
  );
  sg13g2_nor2b_1 _09811_ (
    .A(addr_i_4_),
    .B_N(addr_i_3_),
    .Y(_02645_)
  );
  sg13g2_nand2_1 _09812_ (
    .A(addr_i_2_),
    .B(_02645_),
    .Y(_02656_)
  );
  sg13g2_nand3_1 _09813_ (
    .A(_02623_),
    .B(_02634_),
    .C(_02656_),
    .Y(_02667_)
  );
  sg13g2_o21ai_1 _09814_ (
    .A1(_02613_),
    .A2(_02667_),
    .B1(addr_i_8_),
    .Y(_02678_)
  );
  sg13g2_a22oi_1 _09815_ (
    .A1(_02415_),
    .A2(_02492_),
    .B1(_02580_),
    .B2(_02678_),
    .Y(_02689_)
  );
  sg13g2_buf_1 _09816_ (
    .A(_00374_),
    .X(_02700_)
  );
  sg13g2_a22oi_1 _09817_ (
    .A1(_01932_),
    .A2(_02316_),
    .B1(_02689_),
    .B2(_02700_),
    .Y(_02711_)
  );
  sg13g2_nand2b_1 _09818_ (
    .A_N(addr_i_4_),
    .B(addr_i_3_),
    .Y(_02722_)
  );
  sg13g2_buf_1 _09819_ (
    .A(_02722_),
    .X(_02733_)
  );
  sg13g2_buf_1 _09820_ (
    .A(_02733_),
    .X(_02744_)
  );
  sg13g2_buf_1 _09821_ (
    .A(_00495_),
    .X(_02755_)
  );
  sg13g2_o21ai_1 _09822_ (
    .A1(_02744_),
    .A2(_02755_),
    .B1(addr_i_6_),
    .Y(_02766_)
  );
  sg13g2_buf_1 _09823_ (
    .A(_06496_),
    .X(_02777_)
  );
  sg13g2_nand3b_1 _09824_ (
    .A_N(addr_i_4_),
    .B(addr_i_2_),
    .C(addr_i_5_),
    .Y(_02788_)
  );
  sg13g2_buf_1 _09825_ (
    .A(_02788_),
    .X(_02799_)
  );
  sg13g2_buf_1 _09826_ (
    .A(_02799_),
    .X(_02810_)
  );
  sg13g2_nand2_1 _09827_ (
    .A(_02777_),
    .B(_02810_),
    .Y(_02821_)
  );
  sg13g2_nand3b_1 _09828_ (
    .A_N(addr_i_5_),
    .B(addr_i_2_),
    .C(addr_i_3_),
    .Y(_02832_)
  );
  sg13g2_nand2_1 _09829_ (
    .A(_00462_),
    .B(_02832_),
    .Y(_02843_)
  );
  sg13g2_nand2_1 _09830_ (
    .A(addr_i_4_),
    .B(_02843_),
    .Y(_02854_)
  );
  sg13g2_nand2b_1 _09831_ (
    .A_N(_02821_),
    .B(_02854_),
    .Y(_02865_)
  );
  sg13g2_nand3b_1 _09832_ (
    .A_N(addr_i_5_),
    .B(addr_i_6_),
    .C(addr_i_4_),
    .Y(_02876_)
  );
  sg13g2_buf_1 _09833_ (
    .A(_02876_),
    .X(_02887_)
  );
  sg13g2_buf_1 _09834_ (
    .A(_02887_),
    .X(_02898_)
  );
  sg13g2_nor2b_1 _09835_ (
    .A(addr_i_6_),
    .B_N(addr_i_2_),
    .Y(_02909_)
  );
  sg13g2_nand2_1 _09836_ (
    .A(_00033_),
    .B(_02909_),
    .Y(_02920_)
  );
  sg13g2_buf_1 _09837_ (
    .A(_02920_),
    .X(_02930_)
  );
  sg13g2_a21oi_1 _09838_ (
    .A1(_02898_),
    .A2(_02930_),
    .B1(addr_i_3_),
    .Y(_02941_)
  );
  sg13g2_nor2_1 _09839_ (
    .A(addr_i_9_),
    .B(_01537_),
    .Y(_02952_)
  );
  sg13g2_nand2_1 _09840_ (
    .A(addr_i_7_),
    .B(_02952_),
    .Y(_02963_)
  );
  sg13g2_a22oi_1 _09841_ (
    .A1(_02766_),
    .A2(_02865_),
    .B1(_02941_),
    .B2(_02963_),
    .Y(_02974_)
  );
  sg13g2_a22oi_1 _09842_ (
    .A1(_01351_),
    .A2(_01812_),
    .B1(_02711_),
    .B2(_02974_),
    .Y(_02985_)
  );
  sg13g2_inv_1 _09843_ (
    .A(addr_i_12_),
    .Y(_02996_)
  );
  sg13g2_o21ai_1 _09844_ (
    .A1(addr_i_10_),
    .A2(_02985_),
    .B1(_02996_),
    .Y(_03007_)
  );
  sg13g2_or2_1 _09845_ (
    .A(_01340_),
    .B(_03007_),
    .X(_03018_)
  );
  sg13g2_inv_1 _09846_ (
    .A(addr_i_11_),
    .Y(_03029_)
  );
  sg13g2_buf_1 _09847_ (
    .A(_03029_),
    .X(_03040_)
  );
  sg13g2_buf_1 _09848_ (
    .A(_03040_),
    .X(_03051_)
  );
  sg13g2_buf_1 _09849_ (
    .A(_00791_),
    .X(_03062_)
  );
  sg13g2_nand2_1 _09850_ (
    .A(addr_i_10_),
    .B(_00374_),
    .Y(_03073_)
  );
  sg13g2_nor2_1 _09851_ (
    .A(_03062_),
    .B(_03073_),
    .Y(_03084_)
  );
  sg13g2_and2_1 _09852_ (
    .A(addr_i_4_),
    .B(addr_i_6_),
    .X(_03095_)
  );
  sg13g2_buf_1 _09853_ (
    .A(_03095_),
    .X(_03106_)
  );
  sg13g2_nor2_1 _09854_ (
    .A(addr_i_5_),
    .B(_03106_),
    .Y(_03117_)
  );
  sg13g2_nor2_1 _09855_ (
    .A(addr_i_4_),
    .B(addr_i_6_),
    .Y(_03128_)
  );
  sg13g2_buf_1 _09856_ (
    .A(_03128_),
    .X(_03139_)
  );
  sg13g2_buf_1 _09857_ (
    .A(_03139_),
    .X(_03150_)
  );
  sg13g2_a21oi_1 _09858_ (
    .A1(addr_i_3_),
    .A2(_03117_),
    .B1(_03150_),
    .Y(_03161_)
  );
  sg13g2_buf_1 _09859_ (
    .A(_00539_),
    .X(_03172_)
  );
  sg13g2_and2_1 _09860_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .X(_03183_)
  );
  sg13g2_buf_1 _09861_ (
    .A(_03183_),
    .X(_03194_)
  );
  sg13g2_nand2_1 _09862_ (
    .A(_03172_),
    .B(_03194_),
    .Y(_03205_)
  );
  sg13g2_o21ai_1 _09863_ (
    .A1(addr_i_2_),
    .A2(_03161_),
    .B1(_03205_),
    .Y(_03216_)
  );
  sg13g2_buf_1 _09864_ (
    .A(_01011_),
    .X(_03227_)
  );
  sg13g2_buf_1 _09865_ (
    .A(_03227_),
    .X(_03238_)
  );
  sg13g2_nand2_1 _09866_ (
    .A(addr_i_5_),
    .B(_03238_),
    .Y(_03249_)
  );
  sg13g2_buf_1 _09867_ (
    .A(_01559_),
    .X(_03259_)
  );
  sg13g2_buf_1 _09868_ (
    .A(_07381_),
    .X(_03270_)
  );
  sg13g2_buf_1 _09869_ (
    .A(_03270_),
    .X(_03281_)
  );
  sg13g2_buf_1 _09870_ (
    .A(_03281_),
    .X(_03292_)
  );
  sg13g2_or2_1 _09871_ (
    .A(addr_i_4_),
    .B(addr_i_6_),
    .X(_03303_)
  );
  sg13g2_buf_1 _09872_ (
    .A(_03303_),
    .X(_03314_)
  );
  sg13g2_o21ai_1 _09873_ (
    .A1(addr_i_6_),
    .A2(addr_i_5_),
    .B1(addr_i_4_),
    .Y(_03325_)
  );
  sg13g2_nand2_1 _09874_ (
    .A(_03314_),
    .B(_03325_),
    .Y(_03336_)
  );
  sg13g2_nand2_1 _09875_ (
    .A(addr_i_3_),
    .B(addr_i_7_),
    .Y(_03347_)
  );
  sg13g2_buf_1 _09876_ (
    .A(_03347_),
    .X(_03358_)
  );
  sg13g2_nor2b_1 _09877_ (
    .A(addr_i_3_),
    .B_N(addr_i_4_),
    .Y(_03369_)
  );
  sg13g2_buf_1 _09878_ (
    .A(_03369_),
    .X(_03380_)
  );
  sg13g2_nand2_1 _09879_ (
    .A(_03380_),
    .B(_00550_),
    .Y(_03391_)
  );
  sg13g2_o21ai_1 _09880_ (
    .A1(_03336_),
    .A2(_03358_),
    .B1(_03391_),
    .Y(_03402_)
  );
  sg13g2_nand2_1 _09881_ (
    .A(addr_i_2_),
    .B(addr_i_7_),
    .Y(_03413_)
  );
  sg13g2_buf_1 _09882_ (
    .A(_03413_),
    .X(_03424_)
  );
  sg13g2_inv_1 _09883_ (
    .A(addr_i_5_),
    .Y(_03435_)
  );
  sg13g2_buf_1 _09884_ (
    .A(_03435_),
    .X(_03446_)
  );
  sg13g2_nand2_1 _09885_ (
    .A(_03446_),
    .B(_01439_),
    .Y(_03457_)
  );
  sg13g2_a21oi_1 _09886_ (
    .A1(addr_i_4_),
    .A2(_03424_),
    .B1(_03457_),
    .Y(_03468_)
  );
  sg13g2_or2_1 _09887_ (
    .A(addr_i_2_),
    .B(addr_i_6_),
    .X(_03479_)
  );
  sg13g2_buf_1 _09888_ (
    .A(_03479_),
    .X(_03490_)
  );
  sg13g2_nor2_1 _09889_ (
    .A(addr_i_4_),
    .B(_03490_),
    .Y(_03501_)
  );
  sg13g2_and3_1 _09890_ (
    .A(addr_i_4_),
    .B(addr_i_6_),
    .C(addr_i_5_),
    .X(_03512_)
  );
  sg13g2_buf_1 _09891_ (
    .A(_03512_),
    .X(_03523_)
  );
  sg13g2_nor2_1 _09892_ (
    .A(_03501_),
    .B(_03523_),
    .Y(_03534_)
  );
  sg13g2_o21ai_1 _09893_ (
    .A1(addr_i_2_),
    .A2(addr_i_6_),
    .B1(addr_i_5_),
    .Y(_03545_)
  );
  sg13g2_nor2_1 _09894_ (
    .A(addr_i_4_),
    .B(_03545_),
    .Y(_03555_)
  );
  sg13g2_nor2_1 _09895_ (
    .A(_07933_),
    .B(_01055_),
    .Y(_03566_)
  );
  sg13g2_buf_1 _09896_ (
    .A(_03566_),
    .X(_03577_)
  );
  sg13g2_nor3_1 _09897_ (
    .A(addr_i_3_),
    .B(_03555_),
    .C(_03577_),
    .Y(_03588_)
  );
  sg13g2_a22oi_1 _09898_ (
    .A1(addr_i_3_),
    .A2(_03534_),
    .B1(_03588_),
    .B2(addr_i_7_),
    .Y(_03599_)
  );
  sg13g2_a22oi_1 _09899_ (
    .A1(_03292_),
    .A2(_03402_),
    .B1(_03468_),
    .B2(_03599_),
    .Y(_03610_)
  );
  sg13g2_nor3_1 _09900_ (
    .A(addr_i_4_),
    .B(addr_i_6_),
    .C(addr_i_5_),
    .Y(_03621_)
  );
  sg13g2_buf_1 _09901_ (
    .A(_03621_),
    .X(_03632_)
  );
  sg13g2_nor2_1 _09902_ (
    .A(addr_i_7_),
    .B(_04616_),
    .Y(_03643_)
  );
  sg13g2_nor2_1 _09903_ (
    .A(_03632_),
    .B(_03643_),
    .Y(_03654_)
  );
  sg13g2_buf_1 _09904_ (
    .A(_02645_),
    .X(_03665_)
  );
  sg13g2_buf_1 _09905_ (
    .A(_02097_),
    .X(_03676_)
  );
  sg13g2_nand2_1 _09906_ (
    .A(_03665_),
    .B(_03676_),
    .Y(_03687_)
  );
  sg13g2_o21ai_1 _09907_ (
    .A1(addr_i_3_),
    .A2(_03654_),
    .B1(_03687_),
    .Y(_03698_)
  );
  sg13g2_nand2b_1 _09908_ (
    .A_N(addr_i_6_),
    .B(addr_i_4_),
    .Y(_03709_)
  );
  sg13g2_nor2_1 _09909_ (
    .A(addr_i_3_),
    .B(_03709_),
    .Y(_03720_)
  );
  sg13g2_or2_1 _09910_ (
    .A(addr_i_3_),
    .B(addr_i_6_),
    .X(_03732_)
  );
  sg13g2_buf_1 _09911_ (
    .A(_03732_),
    .X(_03743_)
  );
  sg13g2_o21ai_1 _09912_ (
    .A1(addr_i_4_),
    .A2(addr_i_6_),
    .B1(addr_i_3_),
    .Y(_03754_)
  );
  sg13g2_buf_1 _09913_ (
    .A(_03435_),
    .X(_03765_)
  );
  sg13g2_buf_1 _09914_ (
    .A(_03765_),
    .X(_03776_)
  );
  sg13g2_a21oi_1 _09915_ (
    .A1(_03743_),
    .A2(_03754_),
    .B1(_03776_),
    .Y(_03787_)
  );
  sg13g2_buf_1 _09916_ (
    .A(_00176_),
    .X(_03798_)
  );
  sg13g2_buf_1 _09917_ (
    .A(_03798_),
    .X(_03809_)
  );
  sg13g2_buf_1 _09918_ (
    .A(_03809_),
    .X(_03820_)
  );
  sg13g2_o21ai_1 _09919_ (
    .A1(_03720_),
    .A2(_03787_),
    .B1(_03820_),
    .Y(_03830_)
  );
  sg13g2_nor2_1 _09920_ (
    .A(addr_i_4_),
    .B(addr_i_5_),
    .Y(_03842_)
  );
  sg13g2_buf_1 _09921_ (
    .A(_03842_),
    .X(_03853_)
  );
  sg13g2_nand2b_1 _09922_ (
    .A_N(addr_i_6_),
    .B(addr_i_3_),
    .Y(_03864_)
  );
  sg13g2_nand2b_1 _09923_ (
    .A_N(addr_i_3_),
    .B(addr_i_6_),
    .Y(_03875_)
  );
  sg13g2_nand2_1 _09924_ (
    .A(_03864_),
    .B(_03875_),
    .Y(_03886_)
  );
  sg13g2_nand2_1 _09925_ (
    .A(_03853_),
    .B(_03886_),
    .Y(_03897_)
  );
  sg13g2_buf_1 _09926_ (
    .A(_07381_),
    .X(_03908_)
  );
  sg13g2_buf_1 _09927_ (
    .A(_03908_),
    .X(_03919_)
  );
  sg13g2_buf_1 _09928_ (
    .A(_03919_),
    .X(_03930_)
  );
  sg13g2_a21oi_1 _09929_ (
    .A1(_03830_),
    .A2(_03897_),
    .B1(_03930_),
    .Y(_03941_)
  );
  sg13g2_buf_1 _09930_ (
    .A(_07602_),
    .X(_03953_)
  );
  sg13g2_buf_1 _09931_ (
    .A(_03953_),
    .X(_03964_)
  );
  sg13g2_nand2_1 _09932_ (
    .A(addr_i_8_),
    .B(_03964_),
    .Y(_03975_)
  );
  sg13g2_a22oi_1 _09933_ (
    .A1(_03292_),
    .A2(_03698_),
    .B1(_03941_),
    .B2(_03975_),
    .Y(_03986_)
  );
  sg13g2_a22oi_1 _09934_ (
    .A1(_03259_),
    .A2(_03610_),
    .B1(_03986_),
    .B2(addr_i_9_),
    .Y(_03997_)
  );
  sg13g2_a22oi_1 _09935_ (
    .A1(addr_i_9_),
    .A2(_03249_),
    .B1(_03997_),
    .B2(addr_i_10_),
    .Y(_04008_)
  );
  sg13g2_a22oi_1 _09936_ (
    .A1(_03084_),
    .A2(_03216_),
    .B1(_02996_),
    .B2(_04008_),
    .Y(_04019_)
  );
  sg13g2_nor2_1 _09937_ (
    .A(_03051_),
    .B(_04019_),
    .Y(_04030_)
  );
  sg13g2_buf_1 _09938_ (
    .A(_06496_),
    .X(_04041_)
  );
  sg13g2_buf_1 _09939_ (
    .A(_04041_),
    .X(_04052_)
  );
  sg13g2_nand2b_1 _09940_ (
    .A_N(addr_i_5_),
    .B(addr_i_2_),
    .Y(_04064_)
  );
  sg13g2_buf_1 _09941_ (
    .A(_04064_),
    .X(_04075_)
  );
  sg13g2_buf_1 _09942_ (
    .A(_07159_),
    .X(_04086_)
  );
  sg13g2_a21oi_1 _09943_ (
    .A1(addr_i_3_),
    .A2(_04075_),
    .B1(_04086_),
    .Y(_04097_)
  );
  sg13g2_buf_1 _09944_ (
    .A(_00637_),
    .X(_04108_)
  );
  sg13g2_buf_1 _09945_ (
    .A(_05943_),
    .X(_04119_)
  );
  sg13g2_o21ai_1 _09946_ (
    .A1(_04108_),
    .A2(_04119_),
    .B1(_00297_),
    .Y(_04129_)
  );
  sg13g2_o21ai_1 _09947_ (
    .A1(_09492_),
    .A2(_04097_),
    .B1(_04129_),
    .Y(_04140_)
  );
  sg13g2_buf_1 _09948_ (
    .A(_03369_),
    .X(_04151_)
  );
  sg13g2_buf_1 _09949_ (
    .A(_01373_),
    .X(_04162_)
  );
  sg13g2_nand3_1 _09950_ (
    .A(addr_i_7_),
    .B(_04151_),
    .C(_04162_),
    .Y(_04174_)
  );
  sg13g2_or2_1 _09951_ (
    .A(addr_i_7_),
    .B(addr_i_5_),
    .X(_04185_)
  );
  sg13g2_nor2_1 _09952_ (
    .A(addr_i_2_),
    .B(_04185_),
    .Y(_04196_)
  );
  sg13g2_o21ai_1 _09953_ (
    .A1(_05169_),
    .A2(_04196_),
    .B1(addr_i_3_),
    .Y(_04207_)
  );
  sg13g2_nor2b_1 _09954_ (
    .A(addr_i_3_),
    .B_N(addr_i_2_),
    .Y(_04218_)
  );
  sg13g2_nand2_1 _09955_ (
    .A(_05722_),
    .B(_04218_),
    .Y(_04229_)
  );
  sg13g2_a21o_1 _09956_ (
    .A1(_04207_),
    .A2(_04229_),
    .B1(addr_i_4_),
    .X(_04240_)
  );
  sg13g2_buf_1 _09957_ (
    .A(_00484_),
    .X(_04251_)
  );
  sg13g2_a21oi_1 _09958_ (
    .A1(_04174_),
    .A2(_04240_),
    .B1(_04251_),
    .Y(_04262_)
  );
  sg13g2_a21oi_1 _09959_ (
    .A1(_04052_),
    .A2(_04140_),
    .B1(_04262_),
    .Y(_04273_)
  );
  sg13g2_or3_1 _09960_ (
    .A(addr_i_2_),
    .B(addr_i_7_),
    .C(addr_i_5_),
    .X(_04285_)
  );
  sg13g2_buf_1 _09961_ (
    .A(_04285_),
    .X(_04296_)
  );
  sg13g2_and3_1 _09962_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .C(addr_i_7_),
    .X(_04307_)
  );
  sg13g2_buf_1 _09963_ (
    .A(_04064_),
    .X(_04318_)
  );
  sg13g2_a21oi_1 _09964_ (
    .A1(_04318_),
    .A2(_02338_),
    .B1(addr_i_4_),
    .Y(_04329_)
  );
  sg13g2_o21ai_1 _09965_ (
    .A1(_04307_),
    .A2(_04329_),
    .B1(addr_i_3_),
    .Y(_04340_)
  );
  sg13g2_nand2_1 _09966_ (
    .A(_04296_),
    .B(_04340_),
    .Y(_04351_)
  );
  sg13g2_buf_1 _09967_ (
    .A(_00033_),
    .X(_04362_)
  );
  sg13g2_buf_1 _09968_ (
    .A(_04362_),
    .X(_04373_)
  );
  sg13g2_buf_1 _09969_ (
    .A(_04185_),
    .X(_04384_)
  );
  sg13g2_nand2_1 _09970_ (
    .A(addr_i_2_),
    .B(_01856_),
    .Y(_04396_)
  );
  sg13g2_nand2_1 _09971_ (
    .A(_04384_),
    .B(_04396_),
    .Y(_04407_)
  );
  sg13g2_buf_1 _09972_ (
    .A(_00923_),
    .X(_04418_)
  );
  sg13g2_nand2_1 _09973_ (
    .A(addr_i_4_),
    .B(addr_i_7_),
    .Y(_04429_)
  );
  sg13g2_nor2_1 _09974_ (
    .A(_04418_),
    .B(_04429_),
    .Y(_04439_)
  );
  sg13g2_buf_1 _09975_ (
    .A(_07049_),
    .X(_04450_)
  );
  sg13g2_buf_1 _09976_ (
    .A(_04450_),
    .X(_04461_)
  );
  sg13g2_a22oi_1 _09977_ (
    .A1(_04373_),
    .A2(_04407_),
    .B1(_04439_),
    .B2(_04461_),
    .Y(_04472_)
  );
  sg13g2_nor2_1 _09978_ (
    .A(_00033_),
    .B(_04185_),
    .Y(_04483_)
  );
  sg13g2_nand2b_1 _09979_ (
    .A_N(addr_i_4_),
    .B(addr_i_7_),
    .Y(_04494_)
  );
  sg13g2_nor2_1 _09980_ (
    .A(_00923_),
    .B(_04494_),
    .Y(_04506_)
  );
  sg13g2_or2_1 _09981_ (
    .A(_04483_),
    .B(_04506_),
    .X(_04517_)
  );
  sg13g2_buf_1 _09982_ (
    .A(_01461_),
    .X(_04528_)
  );
  sg13g2_buf_1 _09983_ (
    .A(_04528_),
    .X(_04539_)
  );
  sg13g2_buf_1 _09984_ (
    .A(_03435_),
    .X(_04550_)
  );
  sg13g2_nand2_1 _09985_ (
    .A(addr_i_7_),
    .B(addr_i_6_),
    .Y(_04561_)
  );
  sg13g2_o21ai_1 _09986_ (
    .A1(_04550_),
    .A2(_02547_),
    .B1(_04561_),
    .Y(_04572_)
  );
  sg13g2_a221oi_1 _09987_ (
    .A1(addr_i_2_),
    .A2(_04517_),
    .B1(_04539_),
    .B2(_04572_),
    .C1(addr_i_3_),
    .Y(_04583_)
  );
  sg13g2_nor2_1 _09988_ (
    .A(_04472_),
    .B(_04583_),
    .Y(_04594_)
  );
  sg13g2_a22oi_1 _09989_ (
    .A1(addr_i_6_),
    .A2(_04351_),
    .B1(_04594_),
    .B2(addr_i_8_),
    .Y(_04605_)
  );
  sg13g2_a22oi_1 _09990_ (
    .A1(addr_i_8_),
    .A2(_04273_),
    .B1(_04605_),
    .B2(addr_i_9_),
    .Y(_04617_)
  );
  sg13g2_nand3b_1 _09991_ (
    .A_N(addr_i_2_),
    .B(addr_i_5_),
    .C(addr_i_4_),
    .Y(_04628_)
  );
  sg13g2_a21o_1 _09992_ (
    .A1(_04318_),
    .A2(_04628_),
    .B1(addr_i_3_),
    .X(_04639_)
  );
  sg13g2_nor2b_1 _09993_ (
    .A(addr_i_8_),
    .B_N(addr_i_7_),
    .Y(_04650_)
  );
  sg13g2_nand2_1 _09994_ (
    .A(_06496_),
    .B(_04650_),
    .Y(_04661_)
  );
  sg13g2_buf_1 _09995_ (
    .A(_04661_),
    .X(_04672_)
  );
  sg13g2_nor2_1 _09996_ (
    .A(addr_i_4_),
    .B(_00725_),
    .Y(_04683_)
  );
  sg13g2_nor2_1 _09997_ (
    .A(_04672_),
    .B(_04683_),
    .Y(_04694_)
  );
  sg13g2_buf_1 _09998_ (
    .A(_00385_),
    .X(_04705_)
  );
  sg13g2_nand3_1 _09999_ (
    .A(addr_i_2_),
    .B(addr_i_6_),
    .C(addr_i_5_),
    .Y(_04715_)
  );
  sg13g2_nand2_1 _10000_ (
    .A(_00198_),
    .B(_04715_),
    .Y(_04727_)
  );
  sg13g2_and2_1 _10001_ (
    .A(addr_i_2_),
    .B(addr_i_6_),
    .X(_04738_)
  );
  sg13g2_buf_1 _10002_ (
    .A(_04738_),
    .X(_04749_)
  );
  sg13g2_o21ai_1 _10003_ (
    .A1(_00231_),
    .A2(_04749_),
    .B1(addr_i_7_),
    .Y(_04760_)
  );
  sg13g2_o21ai_1 _10004_ (
    .A1(addr_i_7_),
    .A2(_04727_),
    .B1(_04760_),
    .Y(_04771_)
  );
  sg13g2_nor2_1 _10005_ (
    .A(addr_i_2_),
    .B(_07602_),
    .Y(_04782_)
  );
  sg13g2_buf_1 _10006_ (
    .A(_00912_),
    .X(_04793_)
  );
  sg13g2_nand2b_1 _10007_ (
    .A_N(addr_i_7_),
    .B(addr_i_2_),
    .Y(_04804_)
  );
  sg13g2_nor2_1 _10008_ (
    .A(_04793_),
    .B(_04804_),
    .Y(_04815_)
  );
  sg13g2_o21ai_1 _10009_ (
    .A1(_04782_),
    .A2(_04815_),
    .B1(addr_i_4_),
    .Y(_04826_)
  );
  sg13g2_o21ai_1 _10010_ (
    .A1(addr_i_4_),
    .A2(_04771_),
    .B1(_04826_),
    .Y(_04838_)
  );
  sg13g2_and3_1 _10011_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .C(addr_i_6_),
    .X(_04849_)
  );
  sg13g2_buf_1 _10012_ (
    .A(_00231_),
    .X(_04860_)
  );
  sg13g2_nor3_1 _10013_ (
    .A(addr_i_4_),
    .B(_04860_),
    .C(_04749_),
    .Y(_04871_)
  );
  sg13g2_o21ai_1 _10014_ (
    .A1(_04849_),
    .A2(_04871_),
    .B1(_02053_),
    .Y(_04882_)
  );
  sg13g2_nand2_1 _10015_ (
    .A(addr_i_7_),
    .B(_00231_),
    .Y(_04893_)
  );
  sg13g2_nand2b_1 _10016_ (
    .A_N(addr_i_6_),
    .B(addr_i_7_),
    .Y(_04904_)
  );
  sg13g2_nor2_1 _10017_ (
    .A(_07381_),
    .B(_04904_),
    .Y(_04915_)
  );
  sg13g2_nor2b_1 _10018_ (
    .A(addr_i_7_),
    .B_N(addr_i_2_),
    .Y(_04926_)
  );
  sg13g2_nor2b_1 _10019_ (
    .A(addr_i_2_),
    .B_N(addr_i_6_),
    .Y(_04937_)
  );
  sg13g2_nor3_1 _10020_ (
    .A(addr_i_5_),
    .B(_04926_),
    .C(_04937_),
    .Y(_04949_)
  );
  sg13g2_o21ai_1 _10021_ (
    .A1(_04915_),
    .A2(_04949_),
    .B1(addr_i_4_),
    .Y(_04960_)
  );
  sg13g2_nand3_1 _10022_ (
    .A(_04882_),
    .B(_04893_),
    .C(_04960_),
    .Y(_04971_)
  );
  sg13g2_buf_1 _10023_ (
    .A(_04450_),
    .X(_04981_)
  );
  sg13g2_mux2_1 _10024_ (
    .A0(_04838_),
    .A1(_04971_),
    .S(_04981_),
    .X(_04992_)
  );
  sg13g2_nand2_1 _10025_ (
    .A(_03908_),
    .B(_01636_),
    .Y(_05003_)
  );
  sg13g2_and2_1 _10026_ (
    .A(addr_i_4_),
    .B(addr_i_7_),
    .X(_05014_)
  );
  sg13g2_buf_1 _10027_ (
    .A(_05014_),
    .X(_05025_)
  );
  sg13g2_buf_1 _10028_ (
    .A(_00714_),
    .X(_05036_)
  );
  sg13g2_nand3_1 _10029_ (
    .A(addr_i_3_),
    .B(_05025_),
    .C(_05036_),
    .Y(_05047_)
  );
  sg13g2_o21ai_1 _10030_ (
    .A1(addr_i_3_),
    .A2(_05003_),
    .B1(_05047_),
    .Y(_05059_)
  );
  sg13g2_buf_1 _10031_ (
    .A(_03798_),
    .X(_05070_)
  );
  sg13g2_o21ai_1 _10032_ (
    .A1(addr_i_6_),
    .A2(_02591_),
    .B1(_02009_),
    .Y(_05081_)
  );
  sg13g2_nand2_1 _10033_ (
    .A(addr_i_3_),
    .B(_05081_),
    .Y(_05092_)
  );
  sg13g2_nor2b_1 _10034_ (
    .A(addr_i_6_),
    .B_N(addr_i_3_),
    .Y(_05103_)
  );
  sg13g2_nor2_1 _10035_ (
    .A(addr_i_2_),
    .B(_05103_),
    .Y(_05114_)
  );
  sg13g2_nor2_1 _10036_ (
    .A(addr_i_3_),
    .B(_00231_),
    .Y(_05125_)
  );
  sg13g2_o21ai_1 _10037_ (
    .A1(_05114_),
    .A2(_05125_),
    .B1(addr_i_4_),
    .Y(_05136_)
  );
  sg13g2_and4_1 _10038_ (
    .A(_05070_),
    .B(_05092_),
    .C(_05136_),
    .D(_02799_),
    .X(_05147_)
  );
  sg13g2_a22oi_1 _10039_ (
    .A1(addr_i_6_),
    .A2(_05059_),
    .B1(_05147_),
    .B2(addr_i_8_),
    .Y(_05158_)
  );
  sg13g2_a21oi_1 _10040_ (
    .A1(addr_i_8_),
    .A2(_04992_),
    .B1(_05158_),
    .Y(_05170_)
  );
  sg13g2_a22oi_1 _10041_ (
    .A1(_04639_),
    .A2(_04694_),
    .B1(_04705_),
    .B2(_05170_),
    .Y(_05181_)
  );
  sg13g2_or3_1 _10042_ (
    .A(addr_i_10_),
    .B(_04617_),
    .C(_05181_),
    .X(_05192_)
  );
  sg13g2_nor2_1 _10043_ (
    .A(_03731_),
    .B(_00374_),
    .Y(_05203_)
  );
  sg13g2_buf_1 _10044_ (
    .A(_05203_),
    .X(_05214_)
  );
  sg13g2_buf_1 _10045_ (
    .A(_00066_),
    .X(_05225_)
  );
  sg13g2_buf_1 _10046_ (
    .A(_05225_),
    .X(_05236_)
  );
  sg13g2_buf_1 _10047_ (
    .A(_05236_),
    .X(_05247_)
  );
  sg13g2_buf_1 _10048_ (
    .A(_01153_),
    .X(_05258_)
  );
  sg13g2_buf_1 _10049_ (
    .A(_06938_),
    .X(_05269_)
  );
  sg13g2_buf_1 _10050_ (
    .A(_05269_),
    .X(_05281_)
  );
  sg13g2_nor2_1 _10051_ (
    .A(_05281_),
    .B(_01373_),
    .Y(_05292_)
  );
  sg13g2_buf_1 _10052_ (
    .A(_04362_),
    .X(_05302_)
  );
  sg13g2_o21ai_1 _10053_ (
    .A1(_05258_),
    .A2(_05292_),
    .B1(_05302_),
    .Y(_05313_)
  );
  sg13g2_buf_1 _10054_ (
    .A(_05269_),
    .X(_05324_)
  );
  sg13g2_nor2b_1 _10055_ (
    .A(addr_i_5_),
    .B_N(addr_i_2_),
    .Y(_05335_)
  );
  sg13g2_buf_1 _10056_ (
    .A(_05335_),
    .X(_05346_)
  );
  sg13g2_nand2_1 _10057_ (
    .A(_05324_),
    .B(_05346_),
    .Y(_05357_)
  );
  sg13g2_nand3_1 _10058_ (
    .A(_05247_),
    .B(_05313_),
    .C(_05357_),
    .Y(_05368_)
  );
  sg13g2_buf_1 _10059_ (
    .A(_05103_),
    .X(_05379_)
  );
  sg13g2_nand2_1 _10060_ (
    .A(_01384_),
    .B(_05379_),
    .Y(_05391_)
  );
  sg13g2_buf_1 _10061_ (
    .A(_00637_),
    .X(_05402_)
  );
  sg13g2_a21oi_1 _10062_ (
    .A1(_05357_),
    .A2(_05391_),
    .B1(_05402_),
    .Y(_05413_)
  );
  sg13g2_buf_1 _10063_ (
    .A(_00231_),
    .X(_05424_)
  );
  sg13g2_nand2_1 _10064_ (
    .A(_04218_),
    .B(_05424_),
    .Y(_05435_)
  );
  sg13g2_nand3b_1 _10065_ (
    .A_N(_05413_),
    .B(_05435_),
    .C(addr_i_7_),
    .Y(_05446_)
  );
  sg13g2_buf_1 _10066_ (
    .A(_02031_),
    .X(_05457_)
  );
  sg13g2_a21oi_1 _10067_ (
    .A1(_05457_),
    .A2(_01834_),
    .B1(addr_i_3_),
    .Y(_05468_)
  );
  sg13g2_inv_1 _10068_ (
    .A(_05468_),
    .Y(_05479_)
  );
  sg13g2_nand2_1 _10069_ (
    .A(addr_i_3_),
    .B(_04528_),
    .Y(_05490_)
  );
  sg13g2_nand3_1 _10070_ (
    .A(_01878_),
    .B(_05479_),
    .C(_05490_),
    .Y(_05502_)
  );
  sg13g2_nand4_1 _10071_ (
    .A(addr_i_8_),
    .B(_05368_),
    .C(_05446_),
    .D(_05502_),
    .Y(_05513_)
  );
  sg13g2_buf_1 _10072_ (
    .A(_05390_),
    .X(_05524_)
  );
  sg13g2_nor2_1 _10073_ (
    .A(addr_i_3_),
    .B(_05524_),
    .Y(_05535_)
  );
  sg13g2_buf_1 _10074_ (
    .A(_01899_),
    .X(_05546_)
  );
  sg13g2_nand2_1 _10075_ (
    .A(addr_i_5_),
    .B(_05546_),
    .Y(_05557_)
  );
  sg13g2_buf_1 _10076_ (
    .A(_01910_),
    .X(_05568_)
  );
  sg13g2_nor2_1 _10077_ (
    .A(_02569_),
    .B(_05568_),
    .Y(_05579_)
  );
  sg13g2_o21ai_1 _10078_ (
    .A1(_05535_),
    .A2(_05557_),
    .B1(_05579_),
    .Y(_05589_)
  );
  sg13g2_buf_1 _10079_ (
    .A(_05236_),
    .X(_05600_)
  );
  sg13g2_nand2_1 _10080_ (
    .A(addr_i_5_),
    .B(_02525_),
    .Y(_05612_)
  );
  sg13g2_nand2_1 _10081_ (
    .A(_05600_),
    .B(_05612_),
    .Y(_05623_)
  );
  sg13g2_nor2_1 _10082_ (
    .A(_04550_),
    .B(_04904_),
    .Y(_05634_)
  );
  sg13g2_buf_1 _10083_ (
    .A(_05634_),
    .X(_05645_)
  );
  sg13g2_a21oi_1 _10084_ (
    .A1(_02656_),
    .A2(_05645_),
    .B1(addr_i_8_),
    .Y(_05656_)
  );
  sg13g2_or2_1 _10085_ (
    .A(addr_i_4_),
    .B(addr_i_5_),
    .X(_05667_)
  );
  sg13g2_buf_1 _10086_ (
    .A(_05667_),
    .X(_05678_)
  );
  sg13g2_buf_1 _10087_ (
    .A(_05678_),
    .X(_05689_)
  );
  sg13g2_buf_1 _10088_ (
    .A(_05269_),
    .X(_05700_)
  );
  sg13g2_buf_1 _10089_ (
    .A(_05700_),
    .X(_05711_)
  );
  sg13g2_a21oi_1 _10090_ (
    .A1(_01768_),
    .A2(_05689_),
    .B1(_05711_),
    .Y(_05723_)
  );
  sg13g2_nand2b_1 _10091_ (
    .A_N(addr_i_3_),
    .B(addr_i_4_),
    .Y(_05734_)
  );
  sg13g2_buf_1 _10092_ (
    .A(_05734_),
    .X(_05745_)
  );
  sg13g2_nand2_1 _10093_ (
    .A(addr_i_2_),
    .B(_04793_),
    .Y(_05756_)
  );
  sg13g2_o21ai_1 _10094_ (
    .A1(_05745_),
    .A2(_05756_),
    .B1(_02250_),
    .Y(_05767_)
  );
  sg13g2_o21ai_1 _10095_ (
    .A1(_05723_),
    .A2(_05767_),
    .B1(addr_i_7_),
    .Y(_05778_)
  );
  sg13g2_nand4_1 _10096_ (
    .A(_05589_),
    .B(_05623_),
    .C(_05656_),
    .D(_05778_),
    .Y(_05789_)
  );
  sg13g2_and2_1 _10097_ (
    .A(_05513_),
    .B(_05789_),
    .X(_05800_)
  );
  sg13g2_buf_1 _10098_ (
    .A(_02053_),
    .X(_05811_)
  );
  sg13g2_buf_1 _10099_ (
    .A(_05811_),
    .X(_05822_)
  );
  sg13g2_buf_1 _10100_ (
    .A(_05822_),
    .X(_05834_)
  );
  sg13g2_buf_1 _10101_ (
    .A(_06938_),
    .X(_05845_)
  );
  sg13g2_buf_1 _10102_ (
    .A(_05845_),
    .X(_05856_)
  );
  sg13g2_buf_1 _10103_ (
    .A(_05856_),
    .X(_05867_)
  );
  sg13g2_buf_1 _10104_ (
    .A(_05867_),
    .X(_05877_)
  );
  sg13g2_buf_1 _10105_ (
    .A(_01548_),
    .X(_05888_)
  );
  sg13g2_nand2b_1 _10106_ (
    .A_N(addr_i_4_),
    .B(addr_i_6_),
    .Y(_05899_)
  );
  sg13g2_buf_1 _10107_ (
    .A(_05899_),
    .X(_05910_)
  );
  sg13g2_nand2_1 _10108_ (
    .A(_05546_),
    .B(_05910_),
    .Y(_05921_)
  );
  sg13g2_nor2_1 _10109_ (
    .A(addr_i_5_),
    .B(_01241_),
    .Y(_05932_)
  );
  sg13g2_a21oi_1 _10110_ (
    .A1(addr_i_5_),
    .A2(_05921_),
    .B1(_05932_),
    .Y(_05944_)
  );
  sg13g2_nand2b_1 _10111_ (
    .A_N(addr_i_5_),
    .B(addr_i_8_),
    .Y(_05955_)
  );
  sg13g2_buf_1 _10112_ (
    .A(_00539_),
    .X(_05966_)
  );
  sg13g2_nand2_1 _10113_ (
    .A(_01537_),
    .B(_05966_),
    .Y(_05977_)
  );
  sg13g2_nand2_1 _10114_ (
    .A(_05955_),
    .B(_05977_),
    .Y(_05988_)
  );
  sg13g2_nor2_1 _10115_ (
    .A(_04550_),
    .B(_03709_),
    .Y(_05999_)
  );
  sg13g2_buf_1 _10116_ (
    .A(_05999_),
    .X(_06010_)
  );
  sg13g2_nor2_1 _10117_ (
    .A(_01526_),
    .B(_06386_),
    .Y(_06021_)
  );
  sg13g2_buf_1 _10118_ (
    .A(_02031_),
    .X(_06032_)
  );
  sg13g2_nor3_1 _10119_ (
    .A(addr_i_5_),
    .B(_06021_),
    .C(_06032_),
    .Y(_06043_)
  );
  sg13g2_a22oi_1 _10120_ (
    .A1(addr_i_2_),
    .A2(_05988_),
    .B1(_06010_),
    .B2(_06043_),
    .Y(_06055_)
  );
  sg13g2_o21ai_1 _10121_ (
    .A1(_05888_),
    .A2(_05944_),
    .B1(_06055_),
    .Y(_06066_)
  );
  sg13g2_buf_1 _10122_ (
    .A(_04616_),
    .X(_06077_)
  );
  sg13g2_buf_1 _10123_ (
    .A(_06077_),
    .X(_06088_)
  );
  sg13g2_buf_1 _10124_ (
    .A(_04860_),
    .X(_06099_)
  );
  sg13g2_nand2_1 _10125_ (
    .A(_01548_),
    .B(_06099_),
    .Y(_06110_)
  );
  sg13g2_nand2_1 _10126_ (
    .A(_06088_),
    .B(_06110_),
    .Y(_06121_)
  );
  sg13g2_buf_1 _10127_ (
    .A(_03709_),
    .X(_06132_)
  );
  sg13g2_buf_1 _10128_ (
    .A(_04550_),
    .X(_06143_)
  );
  sg13g2_buf_1 _10129_ (
    .A(_06143_),
    .X(_06154_)
  );
  sg13g2_a22oi_1 _10130_ (
    .A1(addr_i_2_),
    .A2(_06132_),
    .B1(_06154_),
    .B2(addr_i_8_),
    .Y(_06165_)
  );
  sg13g2_buf_1 _10131_ (
    .A(_02909_),
    .X(_06176_)
  );
  sg13g2_nor2b_1 _10132_ (
    .A(addr_i_2_),
    .B_N(addr_i_8_),
    .Y(_06187_)
  );
  sg13g2_buf_1 _10133_ (
    .A(_06187_),
    .X(_06198_)
  );
  sg13g2_nor2b_1 _10134_ (
    .A(addr_i_5_),
    .B_N(addr_i_4_),
    .Y(_06209_)
  );
  sg13g2_buf_1 _10135_ (
    .A(_06209_),
    .X(_06220_)
  );
  sg13g2_o21ai_1 _10136_ (
    .A1(_06176_),
    .A2(_06198_),
    .B1(_06220_),
    .Y(_06231_)
  );
  sg13g2_nand2_1 _10137_ (
    .A(addr_i_3_),
    .B(_06231_),
    .Y(_06242_)
  );
  sg13g2_a22oi_1 _10138_ (
    .A1(_00659_),
    .A2(_06121_),
    .B1(_06165_),
    .B2(_06242_),
    .Y(_06253_)
  );
  sg13g2_nor2_1 _10139_ (
    .A(addr_i_5_),
    .B(_01965_),
    .Y(_06264_)
  );
  sg13g2_buf_1 _10140_ (
    .A(_06264_),
    .X(_06276_)
  );
  sg13g2_a22oi_1 _10141_ (
    .A1(_05877_),
    .A2(_06066_),
    .B1(_06253_),
    .B2(_06276_),
    .Y(_06287_)
  );
  sg13g2_buf_1 _10142_ (
    .A(_05335_),
    .X(_06298_)
  );
  sg13g2_nor2_1 _10143_ (
    .A(_06298_),
    .B(_06198_),
    .Y(_06309_)
  );
  sg13g2_and2_1 _10144_ (
    .A(addr_i_8_),
    .B(addr_i_5_),
    .X(_06320_)
  );
  sg13g2_nor2_1 _10145_ (
    .A(addr_i_2_),
    .B(addr_i_8_),
    .Y(_06331_)
  );
  sg13g2_a21o_1 _10146_ (
    .A1(addr_i_2_),
    .A2(_06320_),
    .B1(_06331_),
    .X(_06342_)
  );
  sg13g2_nor2_1 _10147_ (
    .A(addr_i_3_),
    .B(_06342_),
    .Y(_06353_)
  );
  sg13g2_buf_1 _10148_ (
    .A(_06386_),
    .X(_06364_)
  );
  sg13g2_buf_1 _10149_ (
    .A(_06364_),
    .X(_06375_)
  );
  sg13g2_a22oi_1 _10150_ (
    .A1(addr_i_3_),
    .A2(_06309_),
    .B1(_06353_),
    .B2(_06375_),
    .Y(_06387_)
  );
  sg13g2_buf_1 _10151_ (
    .A(_00539_),
    .X(_06398_)
  );
  sg13g2_nor2b_1 _10152_ (
    .A(addr_i_5_),
    .B_N(addr_i_8_),
    .Y(_06408_)
  );
  sg13g2_buf_1 _10153_ (
    .A(_05281_),
    .X(_06419_)
  );
  sg13g2_a22oi_1 _10154_ (
    .A1(_06398_),
    .A2(_06331_),
    .B1(_06408_),
    .B2(_06419_),
    .Y(_06430_)
  );
  sg13g2_nor2_1 _10155_ (
    .A(addr_i_8_),
    .B(addr_i_5_),
    .Y(_06441_)
  );
  sg13g2_a22oi_1 _10156_ (
    .A1(_06398_),
    .A2(_06198_),
    .B1(_06441_),
    .B2(addr_i_3_),
    .Y(_06452_)
  );
  sg13g2_nor2_1 _10157_ (
    .A(_06430_),
    .B(_06452_),
    .Y(_06463_)
  );
  sg13g2_o21ai_1 _10158_ (
    .A1(_06387_),
    .A2(_06463_),
    .B1(addr_i_4_),
    .Y(_06474_)
  );
  sg13g2_buf_1 _10159_ (
    .A(_02009_),
    .X(_06485_)
  );
  sg13g2_nor2_1 _10160_ (
    .A(_06485_),
    .B(_00813_),
    .Y(_06497_)
  );
  sg13g2_or4_1 _10161_ (
    .A(addr_i_3_),
    .B(addr_i_4_),
    .C(addr_i_2_),
    .D(addr_i_5_),
    .X(_06508_)
  );
  sg13g2_nor2_1 _10162_ (
    .A(_06386_),
    .B(_06508_),
    .Y(_06519_)
  );
  sg13g2_buf_1 _10163_ (
    .A(_00000_),
    .X(_06530_)
  );
  sg13g2_nor3_1 _10164_ (
    .A(addr_i_2_),
    .B(addr_i_6_),
    .C(addr_i_5_),
    .Y(_06541_)
  );
  sg13g2_o21ai_1 _10165_ (
    .A1(_06530_),
    .A2(_06541_),
    .B1(addr_i_3_),
    .Y(_06552_)
  );
  sg13g2_buf_1 _10166_ (
    .A(_04749_),
    .X(_06563_)
  );
  sg13g2_nor3_1 _10167_ (
    .A(addr_i_3_),
    .B(addr_i_2_),
    .C(addr_i_6_),
    .Y(_06574_)
  );
  sg13g2_o21ai_1 _10168_ (
    .A1(_06563_),
    .A2(_06574_),
    .B1(addr_i_5_),
    .Y(_06585_)
  );
  sg13g2_a22oi_1 _10169_ (
    .A1(_06552_),
    .A2(_06585_),
    .B1(addr_i_4_),
    .B2(addr_i_8_),
    .Y(_06596_)
  );
  sg13g2_a22oi_1 _10170_ (
    .A1(addr_i_8_),
    .A2(_06497_),
    .B1(_06519_),
    .B2(_06596_),
    .Y(_06608_)
  );
  sg13g2_buf_1 _10171_ (
    .A(_05070_),
    .X(_06619_)
  );
  sg13g2_buf_1 _10172_ (
    .A(_06619_),
    .X(_06630_)
  );
  sg13g2_a21oi_1 _10173_ (
    .A1(_06474_),
    .A2(_06608_),
    .B1(_06630_),
    .Y(_06641_)
  );
  sg13g2_buf_1 _10174_ (
    .A(_03073_),
    .X(_06652_)
  );
  sg13g2_a22oi_1 _10175_ (
    .A1(_05834_),
    .A2(_06287_),
    .B1(_06641_),
    .B2(_06652_),
    .Y(_06662_)
  );
  sg13g2_a22oi_1 _10176_ (
    .A1(_05214_),
    .A2(_05800_),
    .B1(_02996_),
    .B2(_06662_),
    .Y(_06673_)
  );
  sg13g2_buf_1 _10177_ (
    .A(_01537_),
    .X(_06684_)
  );
  sg13g2_buf_1 _10178_ (
    .A(_06684_),
    .X(_06695_)
  );
  sg13g2_buf_1 _10179_ (
    .A(_06695_),
    .X(_06706_)
  );
  sg13g2_and2_1 _10180_ (
    .A(addr_i_2_),
    .B(addr_i_7_),
    .X(_06718_)
  );
  sg13g2_buf_1 _10181_ (
    .A(_06718_),
    .X(_06729_)
  );
  sg13g2_buf_1 _10182_ (
    .A(_06729_),
    .X(_06740_)
  );
  sg13g2_a22oi_1 _10183_ (
    .A1(addr_i_4_),
    .A2(_01976_),
    .B1(_00890_),
    .B2(addr_i_5_),
    .Y(_06751_)
  );
  sg13g2_or3_1 _10184_ (
    .A(addr_i_3_),
    .B(_06740_),
    .C(_06751_),
    .X(_06762_)
  );
  sg13g2_nand3b_1 _10185_ (
    .A_N(addr_i_6_),
    .B(addr_i_5_),
    .C(addr_i_7_),
    .Y(_06773_)
  );
  sg13g2_buf_1 _10186_ (
    .A(_06773_),
    .X(_06784_)
  );
  sg13g2_buf_1 _10187_ (
    .A(_01153_),
    .X(_06795_)
  );
  sg13g2_buf_1 _10188_ (
    .A(_01033_),
    .X(_06806_)
  );
  sg13g2_o21ai_1 _10189_ (
    .A1(addr_i_7_),
    .A2(_06795_),
    .B1(_06806_),
    .Y(_06817_)
  );
  sg13g2_nand3_1 _10190_ (
    .A(addr_i_3_),
    .B(_06784_),
    .C(_06817_),
    .Y(_06829_)
  );
  sg13g2_nand2b_1 _10191_ (
    .A_N(addr_i_4_),
    .B(addr_i_2_),
    .Y(_06840_)
  );
  sg13g2_buf_1 _10192_ (
    .A(_06840_),
    .X(_06851_)
  );
  sg13g2_buf_1 _10193_ (
    .A(_06851_),
    .X(_06862_)
  );
  sg13g2_buf_1 _10194_ (
    .A(_06862_),
    .X(_06873_)
  );
  sg13g2_buf_1 _10195_ (
    .A(_06485_),
    .X(_06884_)
  );
  sg13g2_buf_1 _10196_ (
    .A(_06884_),
    .X(_06895_)
  );
  sg13g2_buf_1 _10197_ (
    .A(_02064_),
    .X(_06905_)
  );
  sg13g2_a21oi_1 _10198_ (
    .A1(_06873_),
    .A2(_06895_),
    .B1(_06905_),
    .Y(_06916_)
  );
  sg13g2_buf_1 _10199_ (
    .A(_05025_),
    .X(_06927_)
  );
  sg13g2_nor2_1 _10200_ (
    .A(addr_i_4_),
    .B(_04185_),
    .Y(_06939_)
  );
  sg13g2_buf_1 _10201_ (
    .A(_06939_),
    .X(_06950_)
  );
  sg13g2_nor2_1 _10202_ (
    .A(_06927_),
    .B(_06950_),
    .Y(_06961_)
  );
  sg13g2_buf_1 _10203_ (
    .A(_04185_),
    .X(_06972_)
  );
  sg13g2_o21ai_1 _10204_ (
    .A1(_07933_),
    .A2(_06972_),
    .B1(_02591_),
    .Y(_06983_)
  );
  sg13g2_a21oi_1 _10205_ (
    .A1(_06375_),
    .A2(_06983_),
    .B1(addr_i_3_),
    .Y(_06994_)
  );
  sg13g2_a22oi_1 _10206_ (
    .A1(addr_i_3_),
    .A2(_06961_),
    .B1(_06994_),
    .B2(addr_i_2_),
    .Y(_07005_)
  );
  sg13g2_a22oi_1 _10207_ (
    .A1(_06762_),
    .A2(_06829_),
    .B1(_06916_),
    .B2(_07005_),
    .Y(_07016_)
  );
  sg13g2_xor2_1 _10208_ (
    .A(addr_i_7_),
    .B(addr_i_6_),
    .X(_07027_)
  );
  sg13g2_buf_1 _10209_ (
    .A(_07027_),
    .X(_07038_)
  );
  sg13g2_nand2_1 _10210_ (
    .A(addr_i_2_),
    .B(_07038_),
    .Y(_07050_)
  );
  sg13g2_nor2_1 _10211_ (
    .A(addr_i_2_),
    .B(addr_i_7_),
    .Y(_07061_)
  );
  sg13g2_nand2_1 _10212_ (
    .A(addr_i_4_),
    .B(_07061_),
    .Y(_07072_)
  );
  sg13g2_o21ai_1 _10213_ (
    .A1(addr_i_4_),
    .A2(_07050_),
    .B1(_07072_),
    .Y(_07083_)
  );
  sg13g2_nand2_1 _10214_ (
    .A(addr_i_4_),
    .B(_02623_),
    .Y(_07094_)
  );
  sg13g2_buf_1 _10215_ (
    .A(_01856_),
    .X(_07105_)
  );
  sg13g2_nand2_1 _10216_ (
    .A(_07105_),
    .B(_05524_),
    .Y(_07116_)
  );
  sg13g2_nand3_1 _10217_ (
    .A(addr_i_5_),
    .B(_07094_),
    .C(_07116_),
    .Y(_07127_)
  );
  sg13g2_o21ai_1 _10218_ (
    .A1(addr_i_5_),
    .A2(_07083_),
    .B1(_07127_),
    .Y(_07138_)
  );
  sg13g2_buf_1 _10219_ (
    .A(_04981_),
    .X(_07149_)
  );
  sg13g2_buf_1 _10220_ (
    .A(_04561_),
    .X(_07160_)
  );
  sg13g2_nor2_1 _10221_ (
    .A(_04075_),
    .B(_07160_),
    .Y(_07171_)
  );
  sg13g2_nor2_1 _10222_ (
    .A(_07149_),
    .B(_07171_),
    .Y(_07182_)
  );
  sg13g2_nor2_1 _10223_ (
    .A(addr_i_2_),
    .B(_04616_),
    .Y(_07193_)
  );
  sg13g2_o21ai_1 _10224_ (
    .A1(_06176_),
    .A2(_07193_),
    .B1(addr_i_4_),
    .Y(_07204_)
  );
  sg13g2_nor2_1 _10225_ (
    .A(addr_i_2_),
    .B(_04904_),
    .Y(_07215_)
  );
  sg13g2_nor2b_1 _10226_ (
    .A(addr_i_4_),
    .B_N(addr_i_5_),
    .Y(_07226_)
  );
  sg13g2_buf_1 _10227_ (
    .A(_07226_),
    .X(_07237_)
  );
  sg13g2_buf_1 _10228_ (
    .A(_07237_),
    .X(_07248_)
  );
  sg13g2_o21ai_1 _10229_ (
    .A1(_06563_),
    .A2(_07215_),
    .B1(_07248_),
    .Y(_07259_)
  );
  sg13g2_and2_1 _10230_ (
    .A(_07204_),
    .B(_07259_),
    .X(_07271_)
  );
  sg13g2_buf_1 _10231_ (
    .A(_01548_),
    .X(_07282_)
  );
  sg13g2_buf_1 _10232_ (
    .A(_07282_),
    .X(_07293_)
  );
  sg13g2_a221oi_1 _10233_ (
    .A1(_05877_),
    .A2(_07138_),
    .B1(_07182_),
    .B2(_07271_),
    .C1(_07293_),
    .Y(_07304_)
  );
  sg13g2_a21oi_1 _10234_ (
    .A1(_06706_),
    .A2(_07016_),
    .B1(_07304_),
    .Y(_07315_)
  );
  sg13g2_buf_1 _10235_ (
    .A(_00462_),
    .X(_07326_)
  );
  sg13g2_buf_1 _10236_ (
    .A(_07326_),
    .X(_07337_)
  );
  sg13g2_nor2_1 _10237_ (
    .A(addr_i_3_),
    .B(_01241_),
    .Y(_07348_)
  );
  sg13g2_buf_1 _10238_ (
    .A(_01022_),
    .X(_07359_)
  );
  sg13g2_nor2_1 _10239_ (
    .A(_04362_),
    .B(_05346_),
    .Y(_07370_)
  );
  sg13g2_o21ai_1 _10240_ (
    .A1(_07359_),
    .A2(_07370_),
    .B1(addr_i_3_),
    .Y(_07382_)
  );
  sg13g2_nand2b_1 _10241_ (
    .A_N(_07348_),
    .B(_07382_),
    .Y(_07393_)
  );
  sg13g2_buf_1 _10242_ (
    .A(_01494_),
    .X(_07403_)
  );
  sg13g2_a21oi_1 _10243_ (
    .A1(_07337_),
    .A2(_07393_),
    .B1(_07403_),
    .Y(_07414_)
  );
  sg13g2_buf_1 _10244_ (
    .A(_07193_),
    .X(_07425_)
  );
  sg13g2_and2_1 _10245_ (
    .A(addr_i_3_),
    .B(addr_i_4_),
    .X(_07436_)
  );
  sg13g2_buf_1 _10246_ (
    .A(_07436_),
    .X(_07447_)
  );
  sg13g2_buf_1 _10247_ (
    .A(_07447_),
    .X(_07458_)
  );
  sg13g2_nand2b_1 _10248_ (
    .A_N(addr_i_2_),
    .B(addr_i_6_),
    .Y(_07469_)
  );
  sg13g2_o21ai_1 _10249_ (
    .A1(addr_i_5_),
    .A2(_07469_),
    .B1(_00923_),
    .Y(_07480_)
  );
  sg13g2_buf_1 _10250_ (
    .A(_00308_),
    .X(_07492_)
  );
  sg13g2_buf_1 _10251_ (
    .A(_07492_),
    .X(_07503_)
  );
  sg13g2_buf_1 _10252_ (
    .A(_01000_),
    .X(_07514_)
  );
  sg13g2_a221oi_1 _10253_ (
    .A1(_07425_),
    .A2(_07458_),
    .B1(_07480_),
    .B2(_07503_),
    .C1(_07514_),
    .Y(_07525_)
  );
  sg13g2_nand2b_1 _10254_ (
    .A_N(_07525_),
    .B(addr_i_9_),
    .Y(_07536_)
  );
  sg13g2_buf_1 _10255_ (
    .A(_06398_),
    .X(_07547_)
  );
  sg13g2_buf_1 _10256_ (
    .A(_02459_),
    .X(_07558_)
  );
  sg13g2_nand2_1 _10257_ (
    .A(_04450_),
    .B(_05524_),
    .Y(_07569_)
  );
  sg13g2_nand2_1 _10258_ (
    .A(_07558_),
    .B(_07569_),
    .Y(_07580_)
  );
  sg13g2_nand2_1 _10259_ (
    .A(_01526_),
    .B(_03798_),
    .Y(_07591_)
  );
  sg13g2_buf_1 _10260_ (
    .A(_07591_),
    .X(_07603_)
  );
  sg13g2_buf_1 _10261_ (
    .A(_07603_),
    .X(_07614_)
  );
  sg13g2_buf_1 _10262_ (
    .A(_02634_),
    .X(_07625_)
  );
  sg13g2_buf_1 _10263_ (
    .A(_04937_),
    .X(_07636_)
  );
  sg13g2_buf_1 _10264_ (
    .A(_07636_),
    .X(_07647_)
  );
  sg13g2_buf_1 _10265_ (
    .A(_02909_),
    .X(_07658_)
  );
  sg13g2_nor2_1 _10266_ (
    .A(addr_i_3_),
    .B(_07658_),
    .Y(_07668_)
  );
  sg13g2_nor2_1 _10267_ (
    .A(_07647_),
    .B(_07668_),
    .Y(_07679_)
  );
  sg13g2_nor2_1 _10268_ (
    .A(_07625_),
    .B(_07679_),
    .Y(_07690_)
  );
  sg13g2_a22oi_1 _10269_ (
    .A1(_07547_),
    .A2(_07580_),
    .B1(_07614_),
    .B2(_07690_),
    .Y(_07701_)
  );
  sg13g2_nand3b_1 _10270_ (
    .A_N(addr_i_6_),
    .B(addr_i_5_),
    .C(addr_i_4_),
    .Y(_07713_)
  );
  sg13g2_buf_1 _10271_ (
    .A(_07713_),
    .X(_07724_)
  );
  sg13g2_and2_1 _10272_ (
    .A(addr_i_4_),
    .B(addr_i_5_),
    .X(_07735_)
  );
  sg13g2_buf_1 _10273_ (
    .A(_07735_),
    .X(_07746_)
  );
  sg13g2_buf_1 _10274_ (
    .A(_07746_),
    .X(_07757_)
  );
  sg13g2_o21ai_1 _10275_ (
    .A1(_07757_),
    .A2(_03632_),
    .B1(addr_i_3_),
    .Y(_07768_)
  );
  sg13g2_nand2_1 _10276_ (
    .A(_07049_),
    .B(_02108_),
    .Y(_07779_)
  );
  sg13g2_buf_1 _10277_ (
    .A(_07779_),
    .X(_07790_)
  );
  sg13g2_nand3_1 _10278_ (
    .A(_07724_),
    .B(_07768_),
    .C(_07790_),
    .Y(_07801_)
  );
  sg13g2_buf_1 _10279_ (
    .A(_04218_),
    .X(_07812_)
  );
  sg13g2_buf_1 _10280_ (
    .A(_07812_),
    .X(_07824_)
  );
  sg13g2_a221oi_1 _10281_ (
    .A1(_03930_),
    .A2(_07801_),
    .B1(_01044_),
    .B2(_07824_),
    .C1(_00802_),
    .Y(_07835_)
  );
  sg13g2_nor4_1 _10282_ (
    .A(_07414_),
    .B(_07536_),
    .C(_07701_),
    .D(_07835_),
    .Y(_07846_)
  );
  sg13g2_nor2_1 _10283_ (
    .A(_03841_),
    .B(_07846_),
    .Y(_07857_)
  );
  sg13g2_o21ai_1 _10284_ (
    .A1(addr_i_9_),
    .A2(_07315_),
    .B1(_07857_),
    .Y(_07868_)
  );
  sg13g2_buf_1 _10285_ (
    .A(_03842_),
    .X(_07879_)
  );
  sg13g2_buf_1 _10286_ (
    .A(_07879_),
    .X(_07889_)
  );
  sg13g2_xor2_1 _10287_ (
    .A(addr_i_3_),
    .B(addr_i_2_),
    .X(_07900_)
  );
  sg13g2_buf_1 _10288_ (
    .A(_07900_),
    .X(_07911_)
  );
  sg13g2_nor2b_1 _10289_ (
    .A(addr_i_7_),
    .B_N(addr_i_8_),
    .Y(_07922_)
  );
  sg13g2_buf_1 _10290_ (
    .A(_07922_),
    .X(_07934_)
  );
  sg13g2_nand2_1 _10291_ (
    .A(_06607_),
    .B(_07934_),
    .Y(_07945_)
  );
  sg13g2_nor2_1 _10292_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .Y(_07956_)
  );
  sg13g2_buf_1 _10293_ (
    .A(_07956_),
    .X(_07967_)
  );
  sg13g2_nor2_1 _10294_ (
    .A(_07967_),
    .B(_02218_),
    .Y(_07978_)
  );
  sg13g2_a22oi_1 _10295_ (
    .A1(_07889_),
    .A2(_07911_),
    .B1(_07945_),
    .B2(_07978_),
    .Y(_07989_)
  );
  sg13g2_buf_1 _10296_ (
    .A(_03270_),
    .X(_08000_)
  );
  sg13g2_buf_1 _10297_ (
    .A(_08000_),
    .X(_08011_)
  );
  sg13g2_nand2_1 _10298_ (
    .A(_05845_),
    .B(_03842_),
    .Y(_08022_)
  );
  sg13g2_nand2_1 _10299_ (
    .A(_08022_),
    .B(_02207_),
    .Y(_08033_)
  );
  sg13g2_nand2_1 _10300_ (
    .A(addr_i_6_),
    .B(_07922_),
    .Y(_08045_)
  );
  sg13g2_buf_1 _10301_ (
    .A(_07757_),
    .X(_08056_)
  );
  sg13g2_a22oi_1 _10302_ (
    .A1(_08011_),
    .A2(_08033_),
    .B1(_08045_),
    .B2(_08056_),
    .Y(_08067_)
  );
  sg13g2_nor3_1 _10303_ (
    .A(_02700_),
    .B(_07989_),
    .C(_08067_),
    .Y(_08078_)
  );
  sg13g2_nor2b_1 _10304_ (
    .A(addr_i_2_),
    .B_N(addr_i_7_),
    .Y(_08089_)
  );
  sg13g2_buf_1 _10305_ (
    .A(_08089_),
    .X(_08100_)
  );
  sg13g2_buf_1 _10306_ (
    .A(_07447_),
    .X(_08111_)
  );
  sg13g2_nor3_1 _10307_ (
    .A(addr_i_3_),
    .B(addr_i_4_),
    .C(addr_i_7_),
    .Y(_08122_)
  );
  sg13g2_a21oi_1 _10308_ (
    .A1(_08100_),
    .A2(_08111_),
    .B1(_08122_),
    .Y(_08133_)
  );
  sg13g2_buf_1 _10309_ (
    .A(_03194_),
    .X(_08144_)
  );
  sg13g2_buf_1 _10310_ (
    .A(_05269_),
    .X(_08156_)
  );
  sg13g2_buf_1 _10311_ (
    .A(_07226_),
    .X(_08166_)
  );
  sg13g2_nor2_1 _10312_ (
    .A(_08156_),
    .B(_08166_),
    .Y(_08177_)
  );
  sg13g2_buf_1 _10313_ (
    .A(_05225_),
    .X(_08188_)
  );
  sg13g2_o21ai_1 _10314_ (
    .A1(_08144_),
    .A2(_08177_),
    .B1(_08188_),
    .Y(_08199_)
  );
  sg13g2_o21ai_1 _10315_ (
    .A1(_06154_),
    .A2(_08133_),
    .B1(_08199_),
    .Y(_08210_)
  );
  sg13g2_nand3_1 _10316_ (
    .A(addr_i_2_),
    .B(addr_i_7_),
    .C(addr_i_6_),
    .Y(_08221_)
  );
  sg13g2_buf_1 _10317_ (
    .A(_08221_),
    .X(_08232_)
  );
  sg13g2_or2_1 _10318_ (
    .A(addr_i_3_),
    .B(addr_i_5_),
    .X(_08243_)
  );
  sg13g2_buf_1 _10319_ (
    .A(_08243_),
    .X(_08254_)
  );
  sg13g2_buf_1 _10320_ (
    .A(_08254_),
    .X(_08266_)
  );
  sg13g2_a21oi_1 _10321_ (
    .A1(_07072_),
    .A2(_08232_),
    .B1(_08266_),
    .Y(_08277_)
  );
  sg13g2_nor2_1 _10322_ (
    .A(addr_i_2_),
    .B(_02009_),
    .Y(_08288_)
  );
  sg13g2_buf_1 _10323_ (
    .A(_08288_),
    .X(_08299_)
  );
  sg13g2_nor2_1 _10324_ (
    .A(_04904_),
    .B(_00725_),
    .Y(_08310_)
  );
  sg13g2_o21ai_1 _10325_ (
    .A1(_08299_),
    .A2(_08310_),
    .B1(addr_i_3_),
    .Y(_08321_)
  );
  sg13g2_buf_1 _10326_ (
    .A(_02053_),
    .X(_08332_)
  );
  sg13g2_buf_1 _10327_ (
    .A(_04086_),
    .X(_08343_)
  );
  sg13g2_o21ai_1 _10328_ (
    .A1(_08332_),
    .A2(_00616_),
    .B1(_08343_),
    .Y(_08354_)
  );
  sg13g2_a21oi_1 _10329_ (
    .A1(_08321_),
    .A2(_08354_),
    .B1(addr_i_4_),
    .Y(_08365_)
  );
  sg13g2_nor4_1 _10330_ (
    .A(addr_i_8_),
    .B(_08210_),
    .C(_08277_),
    .D(_08365_),
    .Y(_08377_)
  );
  sg13g2_buf_1 _10331_ (
    .A(_08044_),
    .X(_08388_)
  );
  sg13g2_buf_1 _10332_ (
    .A(_08388_),
    .X(_08399_)
  );
  sg13g2_buf_1 _10333_ (
    .A(_07658_),
    .X(_08410_)
  );
  sg13g2_nor2_1 _10334_ (
    .A(_08410_),
    .B(_07425_),
    .Y(_08420_)
  );
  sg13g2_buf_1 _10335_ (
    .A(_01570_),
    .X(_08431_)
  );
  sg13g2_o21ai_1 _10336_ (
    .A1(addr_i_3_),
    .A2(_08420_),
    .B1(_08431_),
    .Y(_08442_)
  );
  sg13g2_nand2_1 _10337_ (
    .A(addr_i_3_),
    .B(addr_i_2_),
    .Y(_08453_)
  );
  sg13g2_buf_1 _10338_ (
    .A(_08453_),
    .X(_08464_)
  );
  sg13g2_nor2_1 _10339_ (
    .A(_06884_),
    .B(_08464_),
    .Y(_08475_)
  );
  sg13g2_buf_1 _10340_ (
    .A(_07514_),
    .X(_08487_)
  );
  sg13g2_a22oi_1 _10341_ (
    .A1(_08399_),
    .A2(_08442_),
    .B1(_08475_),
    .B2(_08487_),
    .Y(_08498_)
  );
  sg13g2_nor2_1 _10342_ (
    .A(_08377_),
    .B(_08498_),
    .Y(_08509_)
  );
  sg13g2_buf_1 _10343_ (
    .A(_03709_),
    .X(_08520_)
  );
  sg13g2_nand2_1 _10344_ (
    .A(addr_i_5_),
    .B(_08520_),
    .Y(_08531_)
  );
  sg13g2_o21ai_1 _10345_ (
    .A1(addr_i_3_),
    .A2(_08531_),
    .B1(_03687_),
    .Y(_08542_)
  );
  sg13g2_buf_1 _10346_ (
    .A(_00835_),
    .X(_08553_)
  );
  sg13g2_buf_1 _10347_ (
    .A(_01899_),
    .X(_08564_)
  );
  sg13g2_nor2_1 _10348_ (
    .A(_09038_),
    .B(_08564_),
    .Y(_08575_)
  );
  sg13g2_a221oi_1 _10349_ (
    .A1(addr_i_2_),
    .A2(_08542_),
    .B1(_08553_),
    .B2(_08575_),
    .C1(_03227_),
    .Y(_08586_)
  );
  sg13g2_buf_1 _10350_ (
    .A(_07967_),
    .X(_08598_)
  );
  sg13g2_nand2_1 _10351_ (
    .A(_01581_),
    .B(_03743_),
    .Y(_08609_)
  );
  sg13g2_o21ai_1 _10352_ (
    .A1(addr_i_4_),
    .A2(_00583_),
    .B1(addr_i_5_),
    .Y(_08620_)
  );
  sg13g2_nor2_1 _10353_ (
    .A(addr_i_6_),
    .B(_08620_),
    .Y(_08631_)
  );
  sg13g2_a21oi_1 _10354_ (
    .A1(_08598_),
    .A2(_08609_),
    .B1(_08631_),
    .Y(_08642_)
  );
  sg13g2_buf_1 _10355_ (
    .A(_05346_),
    .X(_08653_)
  );
  sg13g2_o21ai_1 _10356_ (
    .A1(_08653_),
    .A2(_02130_),
    .B1(addr_i_4_),
    .Y(_08664_)
  );
  sg13g2_buf_1 _10357_ (
    .A(_01494_),
    .X(_08674_)
  );
  sg13g2_a21oi_1 _10358_ (
    .A1(_08642_),
    .A2(_08664_),
    .B1(_08674_),
    .Y(_08685_)
  );
  sg13g2_buf_1 _10359_ (
    .A(_03765_),
    .X(_08696_)
  );
  sg13g2_buf_1 _10360_ (
    .A(_08696_),
    .X(_08708_)
  );
  sg13g2_o21ai_1 _10361_ (
    .A1(addr_i_2_),
    .A2(addr_i_6_),
    .B1(addr_i_3_),
    .Y(_08719_)
  );
  sg13g2_nand2_1 _10362_ (
    .A(_08708_),
    .B(_08719_),
    .Y(_08730_)
  );
  sg13g2_buf_1 _10363_ (
    .A(_07049_),
    .X(_08741_)
  );
  sg13g2_buf_1 _10364_ (
    .A(_08741_),
    .X(_08752_)
  );
  sg13g2_xor2_1 _10365_ (
    .A(addr_i_2_),
    .B(addr_i_6_),
    .X(_08763_)
  );
  sg13g2_buf_1 _10366_ (
    .A(_08763_),
    .X(_08774_)
  );
  sg13g2_buf_1 _10367_ (
    .A(_05845_),
    .X(_08785_)
  );
  sg13g2_buf_1 _10368_ (
    .A(_06077_),
    .X(_08796_)
  );
  sg13g2_nor2_1 _10369_ (
    .A(_08785_),
    .B(_08796_),
    .Y(_08807_)
  );
  sg13g2_a21oi_1 _10370_ (
    .A1(_08752_),
    .A2(_08774_),
    .B1(_08807_),
    .Y(_08819_)
  );
  sg13g2_buf_1 _10371_ (
    .A(_00791_),
    .X(_08830_)
  );
  sg13g2_a22oi_1 _10372_ (
    .A1(_08730_),
    .A2(_08819_),
    .B1(addr_i_4_),
    .B2(_08830_),
    .Y(_08841_)
  );
  sg13g2_buf_1 _10373_ (
    .A(_00583_),
    .X(_08852_)
  );
  sg13g2_xnor2_1 _10374_ (
    .A(addr_i_4_),
    .B(addr_i_5_),
    .Y(_08863_)
  );
  sg13g2_nand2_1 _10375_ (
    .A(_08852_),
    .B(_08863_),
    .Y(_08874_)
  );
  sg13g2_nor2_1 _10376_ (
    .A(addr_i_2_),
    .B(addr_i_5_),
    .Y(_08885_)
  );
  sg13g2_buf_1 _10377_ (
    .A(_08885_),
    .X(_08896_)
  );
  sg13g2_a21oi_1 _10378_ (
    .A1(_08896_),
    .A2(_02733_),
    .B1(_00484_),
    .Y(_08907_)
  );
  sg13g2_a21oi_1 _10379_ (
    .A1(_08874_),
    .A2(_08907_),
    .B1(_07603_),
    .Y(_08918_)
  );
  sg13g2_buf_1 _10380_ (
    .A(_04793_),
    .X(_08930_)
  );
  sg13g2_nand2_1 _10381_ (
    .A(addr_i_3_),
    .B(addr_i_4_),
    .Y(_08941_)
  );
  sg13g2_buf_1 _10382_ (
    .A(_08941_),
    .X(_08951_)
  );
  sg13g2_a22oi_1 _10383_ (
    .A1(_08000_),
    .A2(_08930_),
    .B1(_00791_),
    .B2(_08951_),
    .Y(_08962_)
  );
  sg13g2_or3_1 _10384_ (
    .A(addr_i_9_),
    .B(_08918_),
    .C(_08962_),
    .X(_08973_)
  );
  sg13g2_nor4_1 _10385_ (
    .A(_08586_),
    .B(_08685_),
    .C(_08841_),
    .D(_08973_),
    .Y(_08984_)
  );
  sg13g2_a22oi_1 _10386_ (
    .A1(_08078_),
    .A2(_08509_),
    .B1(_08984_),
    .B2(addr_i_10_),
    .Y(_08995_)
  );
  sg13g2_nor2_1 _10387_ (
    .A(addr_i_12_),
    .B(_08995_),
    .Y(_09006_)
  );
  sg13g2_a221oi_1 _10388_ (
    .A1(_05192_),
    .A2(_06673_),
    .B1(_07868_),
    .B2(_09006_),
    .C1(addr_i_11_),
    .Y(_09017_)
  );
  sg13g2_a21o_1 _10389_ (
    .A1(_03018_),
    .A2(_04030_),
    .B1(_09017_),
    .X(data_o_0_)
  );
  sg13g2_nand2_1 _10390_ (
    .A(_04151_),
    .B(_00495_),
    .Y(_09039_)
  );
  sg13g2_buf_1 _10391_ (
    .A(_04173_),
    .X(_09050_)
  );
  sg13g2_buf_1 _10392_ (
    .A(_09050_),
    .X(_09061_)
  );
  sg13g2_and2_1 _10393_ (
    .A(_09061_),
    .B(_02832_),
    .X(_09072_)
  );
  sg13g2_nor2_1 _10394_ (
    .A(addr_i_5_),
    .B(_06840_),
    .Y(_09083_)
  );
  sg13g2_buf_1 _10395_ (
    .A(_09083_),
    .X(_09094_)
  );
  sg13g2_buf_1 _10396_ (
    .A(_04063_),
    .X(_09105_)
  );
  sg13g2_o21ai_1 _10397_ (
    .A1(addr_i_3_),
    .A2(_09094_),
    .B1(_09105_),
    .Y(_09116_)
  );
  sg13g2_buf_1 _10398_ (
    .A(_01680_),
    .X(_09127_)
  );
  sg13g2_buf_1 _10399_ (
    .A(_09127_),
    .X(_09138_)
  );
  sg13g2_a221oi_1 _10400_ (
    .A1(_09039_),
    .A2(_09072_),
    .B1(_09116_),
    .B2(_09138_),
    .C1(addr_i_8_),
    .Y(_09150_)
  );
  sg13g2_a21oi_1 _10401_ (
    .A1(_00044_),
    .A2(_02909_),
    .B1(_04937_),
    .Y(_09161_)
  );
  sg13g2_nor2_1 _10402_ (
    .A(addr_i_3_),
    .B(_09161_),
    .Y(_09172_)
  );
  sg13g2_nor2_1 _10403_ (
    .A(_05324_),
    .B(_01976_),
    .Y(_09183_)
  );
  sg13g2_nor2_1 _10404_ (
    .A(_09172_),
    .B(_09183_),
    .Y(_09194_)
  );
  sg13g2_buf_1 _10405_ (
    .A(_03864_),
    .X(_09205_)
  );
  sg13g2_nor2_1 _10406_ (
    .A(addr_i_5_),
    .B(_07956_),
    .Y(_09215_)
  );
  sg13g2_buf_1 _10407_ (
    .A(_06530_),
    .X(_09226_)
  );
  sg13g2_a21oi_1 _10408_ (
    .A1(_09226_),
    .A2(_00319_),
    .B1(addr_i_7_),
    .Y(_09237_)
  );
  sg13g2_o21ai_1 _10409_ (
    .A1(_09205_),
    .A2(_09215_),
    .B1(_09237_),
    .Y(_09248_)
  );
  sg13g2_buf_1 _10410_ (
    .A(_01406_),
    .X(_09260_)
  );
  sg13g2_buf_1 _10411_ (
    .A(_04108_),
    .X(_09271_)
  );
  sg13g2_a21oi_1 _10412_ (
    .A1(_09260_),
    .A2(_03457_),
    .B1(_09271_),
    .Y(_09282_)
  );
  sg13g2_nor2_1 _10413_ (
    .A(_09248_),
    .B(_09282_),
    .Y(_09293_)
  );
  sg13g2_o21ai_1 _10414_ (
    .A1(addr_i_5_),
    .A2(_09194_),
    .B1(_09293_),
    .Y(_09304_)
  );
  sg13g2_buf_1 _10415_ (
    .A(_00374_),
    .X(_09315_)
  );
  sg13g2_buf_1 _10416_ (
    .A(_09315_),
    .X(_09326_)
  );
  sg13g2_a21oi_1 _10417_ (
    .A1(_09150_),
    .A2(_09304_),
    .B1(_09326_),
    .Y(_09337_)
  );
  sg13g2_nor2_1 _10418_ (
    .A(_07491_),
    .B(_00923_),
    .Y(_09348_)
  );
  sg13g2_buf_1 _10419_ (
    .A(_09348_),
    .X(_09359_)
  );
  sg13g2_buf_1 _10420_ (
    .A(_01055_),
    .X(_09371_)
  );
  sg13g2_nand2_1 _10421_ (
    .A(_08696_),
    .B(_09371_),
    .Y(_09382_)
  );
  sg13g2_buf_1 _10422_ (
    .A(_01965_),
    .X(_09393_)
  );
  sg13g2_or3_1 _10423_ (
    .A(addr_i_2_),
    .B(addr_i_6_),
    .C(addr_i_5_),
    .X(_09404_)
  );
  sg13g2_buf_1 _10424_ (
    .A(_09404_),
    .X(_09415_)
  );
  sg13g2_nand3_1 _10425_ (
    .A(addr_i_3_),
    .B(_09393_),
    .C(_09415_),
    .Y(_09426_)
  );
  sg13g2_o21ai_1 _10426_ (
    .A1(addr_i_3_),
    .A2(_09382_),
    .B1(_09426_),
    .Y(_09437_)
  );
  sg13g2_nand2_1 _10427_ (
    .A(_04318_),
    .B(_04418_),
    .Y(_09448_)
  );
  sg13g2_buf_1 _10428_ (
    .A(_03676_),
    .X(_09459_)
  );
  sg13g2_a22oi_1 _10429_ (
    .A1(addr_i_3_),
    .A2(_09448_),
    .B1(_09459_),
    .B2(addr_i_4_),
    .Y(_09469_)
  );
  sg13g2_a21oi_1 _10430_ (
    .A1(addr_i_4_),
    .A2(_09437_),
    .B1(_09469_),
    .Y(_09471_)
  );
  sg13g2_o21ai_1 _10431_ (
    .A1(_09359_),
    .A2(_09471_),
    .B1(addr_i_7_),
    .Y(_09472_)
  );
  sg13g2_buf_1 _10432_ (
    .A(_07105_),
    .X(_09473_)
  );
  sg13g2_buf_1 _10433_ (
    .A(_09473_),
    .X(_09474_)
  );
  sg13g2_nand2_1 _10434_ (
    .A(_03435_),
    .B(_05390_),
    .Y(_09475_)
  );
  sg13g2_buf_1 _10435_ (
    .A(_09475_),
    .X(_09476_)
  );
  sg13g2_nand2_1 _10436_ (
    .A(_05845_),
    .B(_01142_),
    .Y(_09477_)
  );
  sg13g2_buf_1 _10437_ (
    .A(_09477_),
    .X(_09478_)
  );
  sg13g2_nand2_1 _10438_ (
    .A(addr_i_3_),
    .B(_00736_),
    .Y(_09479_)
  );
  sg13g2_nand3_1 _10439_ (
    .A(addr_i_4_),
    .B(_09478_),
    .C(_09479_),
    .Y(_09480_)
  );
  sg13g2_nand3_1 _10440_ (
    .A(_09474_),
    .B(_09476_),
    .C(_09480_),
    .Y(_09482_)
  );
  sg13g2_nand2_1 _10441_ (
    .A(addr_i_4_),
    .B(_00495_),
    .Y(_09483_)
  );
  sg13g2_and2_1 _10442_ (
    .A(_01087_),
    .B(_09483_),
    .X(_09484_)
  );
  sg13g2_buf_1 _10443_ (
    .A(_05225_),
    .X(_09485_)
  );
  sg13g2_buf_1 _10444_ (
    .A(_09485_),
    .X(_09486_)
  );
  sg13g2_buf_1 _10445_ (
    .A(_09486_),
    .X(_09487_)
  );
  sg13g2_o21ai_1 _10446_ (
    .A1(addr_i_3_),
    .A2(_09484_),
    .B1(_09487_),
    .Y(_09488_)
  );
  sg13g2_nand4_1 _10447_ (
    .A(addr_i_8_),
    .B(_09472_),
    .C(_09482_),
    .D(_09488_),
    .Y(_09489_)
  );
  sg13g2_nand2_1 _10448_ (
    .A(_09337_),
    .B(_09489_),
    .Y(_09490_)
  );
  sg13g2_buf_1 _10449_ (
    .A(_08156_),
    .X(_09491_)
  );
  sg13g2_buf_1 _10450_ (
    .A(_06209_),
    .X(_09493_)
  );
  sg13g2_buf_1 _10451_ (
    .A(_09493_),
    .X(_09494_)
  );
  sg13g2_nor2_1 _10452_ (
    .A(addr_i_4_),
    .B(_02371_),
    .Y(_09495_)
  );
  sg13g2_nor3_1 _10453_ (
    .A(_09491_),
    .B(_09494_),
    .C(_09495_),
    .Y(_09496_)
  );
  sg13g2_buf_1 _10454_ (
    .A(_07746_),
    .X(_09497_)
  );
  sg13g2_nor2_1 _10455_ (
    .A(addr_i_5_),
    .B(_02283_),
    .Y(_09498_)
  );
  sg13g2_buf_1 _10456_ (
    .A(_09498_),
    .X(_09499_)
  );
  sg13g2_nor3_1 _10457_ (
    .A(addr_i_3_),
    .B(_09497_),
    .C(_09499_),
    .Y(_09500_)
  );
  sg13g2_nor2b_1 _10458_ (
    .A(addr_i_7_),
    .B_N(addr_i_4_),
    .Y(_09501_)
  );
  sg13g2_nor2_1 _10459_ (
    .A(addr_i_4_),
    .B(_04904_),
    .Y(_09502_)
  );
  sg13g2_nor2_1 _10460_ (
    .A(_09501_),
    .B(_09502_),
    .Y(_09504_)
  );
  sg13g2_o21ai_1 _10461_ (
    .A1(_09496_),
    .A2(_09500_),
    .B1(_09504_),
    .Y(_09505_)
  );
  sg13g2_and3_1 _10462_ (
    .A(addr_i_7_),
    .B(addr_i_6_),
    .C(addr_i_5_),
    .X(_09506_)
  );
  sg13g2_buf_1 _10463_ (
    .A(_09506_),
    .X(_09507_)
  );
  sg13g2_nand2_1 _10464_ (
    .A(_05281_),
    .B(_02558_),
    .Y(_09508_)
  );
  sg13g2_buf_1 _10465_ (
    .A(_04429_),
    .X(_09509_)
  );
  sg13g2_buf_1 _10466_ (
    .A(_02020_),
    .X(_09510_)
  );
  sg13g2_nand3_1 _10467_ (
    .A(addr_i_3_),
    .B(_09509_),
    .C(_09510_),
    .Y(_09511_)
  );
  sg13g2_o21ai_1 _10468_ (
    .A1(_09507_),
    .A2(_09508_),
    .B1(_09511_),
    .Y(_09512_)
  );
  sg13g2_buf_1 _10469_ (
    .A(_05734_),
    .X(_09513_)
  );
  sg13g2_buf_1 _10470_ (
    .A(_05722_),
    .X(_00001_)
  );
  sg13g2_a22oi_1 _10471_ (
    .A1(addr_i_6_),
    .A2(_09513_),
    .B1(_00001_),
    .B2(_09061_),
    .Y(_00002_)
  );
  sg13g2_nor2_1 _10472_ (
    .A(addr_i_8_),
    .B(_00002_),
    .Y(_00003_)
  );
  sg13g2_o21ai_1 _10473_ (
    .A1(addr_i_2_),
    .A2(_09512_),
    .B1(_00003_),
    .Y(_00004_)
  );
  sg13g2_a21oi_1 _10474_ (
    .A1(addr_i_2_),
    .A2(_09505_),
    .B1(_00004_),
    .Y(_00005_)
  );
  sg13g2_buf_1 _10475_ (
    .A(_04561_),
    .X(_00006_)
  );
  sg13g2_buf_1 _10476_ (
    .A(_00006_),
    .X(_00007_)
  );
  sg13g2_xor2_1 _10477_ (
    .A(addr_i_4_),
    .B(addr_i_5_),
    .X(_00008_)
  );
  sg13g2_nor2_1 _10478_ (
    .A(addr_i_3_),
    .B(_00008_),
    .Y(_00009_)
  );
  sg13g2_buf_1 _10479_ (
    .A(_01856_),
    .X(_00010_)
  );
  sg13g2_nand2_1 _10480_ (
    .A(_00010_),
    .B(_09478_),
    .Y(_00012_)
  );
  sg13g2_o21ai_1 _10481_ (
    .A1(_00007_),
    .A2(_00009_),
    .B1(_00012_),
    .Y(_00013_)
  );
  sg13g2_buf_1 _10482_ (
    .A(_07159_),
    .X(_00014_)
  );
  sg13g2_buf_1 _10483_ (
    .A(_00014_),
    .X(_00015_)
  );
  sg13g2_buf_1 _10484_ (
    .A(_04804_),
    .X(_00016_)
  );
  sg13g2_nor2_1 _10485_ (
    .A(_08044_),
    .B(_00016_),
    .Y(_00017_)
  );
  sg13g2_o21ai_1 _10486_ (
    .A1(_00015_),
    .A2(_00017_),
    .B1(addr_i_3_),
    .Y(_00018_)
  );
  sg13g2_buf_1 _10487_ (
    .A(_00451_),
    .X(_00019_)
  );
  sg13g2_buf_1 _10488_ (
    .A(_00019_),
    .X(_00020_)
  );
  sg13g2_buf_1 _10489_ (
    .A(_02283_),
    .X(_00021_)
  );
  sg13g2_nor2_1 _10490_ (
    .A(_00020_),
    .B(_00021_),
    .Y(_00023_)
  );
  sg13g2_buf_1 _10491_ (
    .A(_04075_),
    .X(_00024_)
  );
  sg13g2_buf_1 _10492_ (
    .A(_04904_),
    .X(_00025_)
  );
  sg13g2_nor2_1 _10493_ (
    .A(_00024_),
    .B(_00025_),
    .Y(_00026_)
  );
  sg13g2_o21ai_1 _10494_ (
    .A1(_09486_),
    .A2(_00026_),
    .B1(addr_i_4_),
    .Y(_00027_)
  );
  sg13g2_nand2b_1 _10495_ (
    .A_N(_00023_),
    .B(_00027_),
    .Y(_00028_)
  );
  sg13g2_buf_1 _10496_ (
    .A(_00209_),
    .X(_00029_)
  );
  sg13g2_buf_1 _10497_ (
    .A(_05734_),
    .X(_00030_)
  );
  sg13g2_nor2_1 _10498_ (
    .A(addr_i_2_),
    .B(_00030_),
    .Y(_00031_)
  );
  sg13g2_buf_1 _10499_ (
    .A(_00025_),
    .X(_00032_)
  );
  sg13g2_buf_1 _10500_ (
    .A(_02722_),
    .X(_00034_)
  );
  sg13g2_nor3_1 _10501_ (
    .A(_08653_),
    .B(_00032_),
    .C(_00034_),
    .Y(_00035_)
  );
  sg13g2_a22oi_1 _10502_ (
    .A1(_00029_),
    .A2(_00031_),
    .B1(_00035_),
    .B2(_05888_),
    .Y(_00036_)
  );
  sg13g2_nand2_1 _10503_ (
    .A(_05324_),
    .B(_05225_),
    .Y(_00037_)
  );
  sg13g2_xor2_1 _10504_ (
    .A(addr_i_2_),
    .B(addr_i_5_),
    .X(_00038_)
  );
  sg13g2_nand2_1 _10505_ (
    .A(addr_i_4_),
    .B(_00038_),
    .Y(_00039_)
  );
  sg13g2_nand2b_1 _10506_ (
    .A_N(_00037_),
    .B(_00039_),
    .Y(_00040_)
  );
  sg13g2_nand2_1 _10507_ (
    .A(_00036_),
    .B(_00040_),
    .Y(_00041_)
  );
  sg13g2_a221oi_1 _10508_ (
    .A1(_00013_),
    .A2(_00018_),
    .B1(_00028_),
    .B2(addr_i_3_),
    .C1(_00041_),
    .Y(_00042_)
  );
  sg13g2_nor3_1 _10509_ (
    .A(addr_i_9_),
    .B(_00005_),
    .C(_00042_),
    .Y(_00043_)
  );
  sg13g2_nor2_1 _10510_ (
    .A(addr_i_10_),
    .B(_00043_),
    .Y(_00045_)
  );
  sg13g2_buf_1 _10511_ (
    .A(_05281_),
    .X(_00046_)
  );
  sg13g2_buf_1 _10512_ (
    .A(_00046_),
    .X(_00047_)
  );
  sg13g2_buf_1 _10513_ (
    .A(_00047_),
    .X(_00048_)
  );
  sg13g2_nand2_1 _10514_ (
    .A(_00176_),
    .B(_00539_),
    .Y(_00049_)
  );
  sg13g2_buf_1 _10515_ (
    .A(_00049_),
    .X(_00050_)
  );
  sg13g2_buf_1 _10516_ (
    .A(_00050_),
    .X(_00051_)
  );
  sg13g2_buf_1 _10517_ (
    .A(_07160_),
    .X(_00052_)
  );
  sg13g2_buf_1 _10518_ (
    .A(_00052_),
    .X(_00053_)
  );
  sg13g2_o21ai_1 _10519_ (
    .A1(_06873_),
    .A2(_00051_),
    .B1(_00053_),
    .Y(_00054_)
  );
  sg13g2_buf_1 _10520_ (
    .A(_04893_),
    .X(_00056_)
  );
  sg13g2_nor2_1 _10521_ (
    .A(addr_i_4_),
    .B(_02283_),
    .Y(_00057_)
  );
  sg13g2_o21ai_1 _10522_ (
    .A1(_06010_),
    .A2(_00057_),
    .B1(addr_i_2_),
    .Y(_00058_)
  );
  sg13g2_buf_1 _10523_ (
    .A(_05700_),
    .X(_00059_)
  );
  sg13g2_buf_1 _10524_ (
    .A(_00059_),
    .X(_00060_)
  );
  sg13g2_buf_1 _10525_ (
    .A(_00060_),
    .X(_00061_)
  );
  sg13g2_a21oi_1 _10526_ (
    .A1(_00056_),
    .A2(_00058_),
    .B1(_00061_),
    .Y(_00062_)
  );
  sg13g2_a21oi_1 _10527_ (
    .A1(_00048_),
    .A2(_00054_),
    .B1(_00062_),
    .Y(_00063_)
  );
  sg13g2_buf_1 _10528_ (
    .A(_07381_),
    .X(_00064_)
  );
  sg13g2_buf_1 _10529_ (
    .A(_00064_),
    .X(_00065_)
  );
  sg13g2_buf_1 _10530_ (
    .A(_00065_),
    .X(_00067_)
  );
  sg13g2_buf_1 _10531_ (
    .A(_00067_),
    .X(_00068_)
  );
  sg13g2_buf_1 _10532_ (
    .A(_06972_),
    .X(_00069_)
  );
  sg13g2_buf_1 _10533_ (
    .A(_04429_),
    .X(_00070_)
  );
  sg13g2_nand3_1 _10534_ (
    .A(addr_i_3_),
    .B(_00069_),
    .C(_00070_),
    .Y(_00071_)
  );
  sg13g2_buf_1 _10535_ (
    .A(_03380_),
    .X(_00072_)
  );
  sg13g2_buf_1 _10536_ (
    .A(_00072_),
    .X(_00073_)
  );
  sg13g2_nand2_1 _10537_ (
    .A(addr_i_5_),
    .B(_02547_),
    .Y(_00074_)
  );
  sg13g2_a21oi_1 _10538_ (
    .A1(_00073_),
    .A2(_00074_),
    .B1(_09495_),
    .Y(_00075_)
  );
  sg13g2_nand2_1 _10539_ (
    .A(_00071_),
    .B(_00075_),
    .Y(_00076_)
  );
  sg13g2_nand2_1 _10540_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .Y(_00078_)
  );
  sg13g2_buf_1 _10541_ (
    .A(_00078_),
    .X(_00079_)
  );
  sg13g2_buf_1 _10542_ (
    .A(_00079_),
    .X(_00080_)
  );
  sg13g2_nor2_1 _10543_ (
    .A(_03964_),
    .B(_00080_),
    .Y(_00081_)
  );
  sg13g2_a22oi_1 _10544_ (
    .A1(_00068_),
    .A2(_00076_),
    .B1(_00081_),
    .B2(addr_i_8_),
    .Y(_00082_)
  );
  sg13g2_buf_1 _10545_ (
    .A(_00956_),
    .X(_00083_)
  );
  sg13g2_buf_1 _10546_ (
    .A(_00083_),
    .X(_00084_)
  );
  sg13g2_nor2_1 _10547_ (
    .A(_05600_),
    .B(_00029_),
    .Y(_00085_)
  );
  sg13g2_buf_1 _10548_ (
    .A(_04926_),
    .X(_00086_)
  );
  sg13g2_nor2_1 _10549_ (
    .A(addr_i_2_),
    .B(_04561_),
    .Y(_00087_)
  );
  sg13g2_o21ai_1 _10550_ (
    .A1(_00086_),
    .A2(_00087_),
    .B1(_06143_),
    .Y(_00089_)
  );
  sg13g2_nor2_1 _10551_ (
    .A(_04550_),
    .B(_04926_),
    .Y(_00090_)
  );
  sg13g2_buf_1 _10552_ (
    .A(_06364_),
    .X(_00091_)
  );
  sg13g2_o21ai_1 _10553_ (
    .A1(_00001_),
    .A2(_00090_),
    .B1(_00091_),
    .Y(_00092_)
  );
  sg13g2_and3_1 _10554_ (
    .A(addr_i_4_),
    .B(_00089_),
    .C(_00092_),
    .X(_00093_)
  );
  sg13g2_a21oi_1 _10555_ (
    .A1(_00084_),
    .A2(_00085_),
    .B1(_00093_),
    .Y(_00094_)
  );
  sg13g2_a21oi_1 _10556_ (
    .A1(addr_i_7_),
    .A2(_01066_),
    .B1(addr_i_4_),
    .Y(_00095_)
  );
  sg13g2_nor2_1 _10557_ (
    .A(addr_i_2_),
    .B(_02558_),
    .Y(_00096_)
  );
  sg13g2_nor2_1 _10558_ (
    .A(_00095_),
    .B(_00096_),
    .Y(_00097_)
  );
  sg13g2_nor2_1 _10559_ (
    .A(_03798_),
    .B(_04937_),
    .Y(_00098_)
  );
  sg13g2_nor2_1 _10560_ (
    .A(_03908_),
    .B(_02558_),
    .Y(_00100_)
  );
  sg13g2_a22oi_1 _10561_ (
    .A1(addr_i_4_),
    .A2(_00098_),
    .B1(_00100_),
    .B2(addr_i_5_),
    .Y(_00101_)
  );
  sg13g2_a22oi_1 _10562_ (
    .A1(addr_i_5_),
    .A2(_00097_),
    .B1(_00101_),
    .B2(addr_i_3_),
    .Y(_00102_)
  );
  sg13g2_buf_1 _10563_ (
    .A(_00016_),
    .X(_00103_)
  );
  sg13g2_buf_1 _10564_ (
    .A(_02591_),
    .X(_00104_)
  );
  sg13g2_buf_1 _10565_ (
    .A(_00104_),
    .X(_00105_)
  );
  sg13g2_o21ai_1 _10566_ (
    .A1(_00103_),
    .A2(_00105_),
    .B1(addr_i_8_),
    .Y(_00106_)
  );
  sg13g2_a22oi_1 _10567_ (
    .A1(addr_i_3_),
    .A2(_00094_),
    .B1(_00102_),
    .B2(_00106_),
    .Y(_00107_)
  );
  sg13g2_nand2_1 _10568_ (
    .A(addr_i_10_),
    .B(addr_i_9_),
    .Y(_00108_)
  );
  sg13g2_buf_1 _10569_ (
    .A(_00108_),
    .X(_00109_)
  );
  sg13g2_a22oi_1 _10570_ (
    .A1(_00063_),
    .A2(_00082_),
    .B1(_00107_),
    .B2(_00109_),
    .Y(_00111_)
  );
  sg13g2_buf_1 _10571_ (
    .A(_01548_),
    .X(_00112_)
  );
  sg13g2_buf_1 _10572_ (
    .A(_00112_),
    .X(_00113_)
  );
  sg13g2_buf_1 _10573_ (
    .A(_00113_),
    .X(_00114_)
  );
  sg13g2_buf_1 _10574_ (
    .A(_02086_),
    .X(_00115_)
  );
  sg13g2_buf_1 _10575_ (
    .A(_00115_),
    .X(_00116_)
  );
  sg13g2_buf_1 _10576_ (
    .A(_04550_),
    .X(_00117_)
  );
  sg13g2_nand2_1 _10577_ (
    .A(_00117_),
    .B(_03314_),
    .Y(_00118_)
  );
  sg13g2_nor2_1 _10578_ (
    .A(addr_i_4_),
    .B(_04616_),
    .Y(_00119_)
  );
  sg13g2_buf_1 _10579_ (
    .A(_07491_),
    .X(_00120_)
  );
  sg13g2_buf_1 _10580_ (
    .A(_00120_),
    .X(_00122_)
  );
  sg13g2_buf_1 _10581_ (
    .A(_00122_),
    .X(_00123_)
  );
  sg13g2_a22oi_1 _10582_ (
    .A1(_00116_),
    .A2(_00118_),
    .B1(_00119_),
    .B2(_00123_),
    .Y(_00124_)
  );
  sg13g2_nand2_1 _10583_ (
    .A(addr_i_4_),
    .B(_04793_),
    .Y(_00125_)
  );
  sg13g2_a21o_1 _10584_ (
    .A1(_05114_),
    .A2(_00125_),
    .B1(addr_i_7_),
    .X(_00126_)
  );
  sg13g2_nor2_1 _10585_ (
    .A(_05700_),
    .B(_02525_),
    .Y(_00127_)
  );
  sg13g2_buf_1 _10586_ (
    .A(_06099_),
    .X(_00128_)
  );
  sg13g2_o21ai_1 _10587_ (
    .A1(_04307_),
    .A2(_00127_),
    .B1(_00128_),
    .Y(_00129_)
  );
  sg13g2_o21ai_1 _10588_ (
    .A1(_00124_),
    .A2(_00126_),
    .B1(_00129_),
    .Y(_00130_)
  );
  sg13g2_nand2_1 _10589_ (
    .A(_05943_),
    .B(_05966_),
    .Y(_00131_)
  );
  sg13g2_a21oi_1 _10590_ (
    .A1(addr_i_4_),
    .A2(_04162_),
    .B1(addr_i_3_),
    .Y(_00133_)
  );
  sg13g2_o21ai_1 _10591_ (
    .A1(_07889_),
    .A2(_00133_),
    .B1(addr_i_6_),
    .Y(_00134_)
  );
  sg13g2_a21oi_1 _10592_ (
    .A1(_00131_),
    .A2(_00134_),
    .B1(_03062_),
    .Y(_00135_)
  );
  sg13g2_nor2_1 _10593_ (
    .A(_06154_),
    .B(_07647_),
    .Y(_00136_)
  );
  sg13g2_nand2_1 _10594_ (
    .A(_07491_),
    .B(_02108_),
    .Y(_00137_)
  );
  sg13g2_buf_1 _10595_ (
    .A(_00137_),
    .X(_00138_)
  );
  sg13g2_o21ai_1 _10596_ (
    .A1(addr_i_3_),
    .A2(_00136_),
    .B1(_00138_),
    .Y(_00139_)
  );
  sg13g2_nand2_1 _10597_ (
    .A(addr_i_3_),
    .B(_02020_),
    .Y(_00140_)
  );
  sg13g2_nor2_1 _10598_ (
    .A(_07824_),
    .B(_00561_),
    .Y(_00141_)
  );
  sg13g2_a21oi_1 _10599_ (
    .A1(_00140_),
    .A2(_00141_),
    .B1(addr_i_4_),
    .Y(_00142_)
  );
  sg13g2_a22oi_1 _10600_ (
    .A1(addr_i_4_),
    .A2(_00139_),
    .B1(_00142_),
    .B2(_09359_),
    .Y(_00144_)
  );
  sg13g2_buf_1 _10601_ (
    .A(_03270_),
    .X(_00145_)
  );
  sg13g2_buf_1 _10602_ (
    .A(_00145_),
    .X(_00146_)
  );
  sg13g2_or3_1 _10603_ (
    .A(addr_i_4_),
    .B(addr_i_6_),
    .C(addr_i_5_),
    .X(_00147_)
  );
  sg13g2_buf_1 _10604_ (
    .A(_00147_),
    .X(_00148_)
  );
  sg13g2_nand2_1 _10605_ (
    .A(_01252_),
    .B(_00148_),
    .Y(_00149_)
  );
  sg13g2_buf_1 _10606_ (
    .A(_01384_),
    .X(_00150_)
  );
  sg13g2_buf_1 _10607_ (
    .A(_03314_),
    .X(_00151_)
  );
  sg13g2_a21oi_1 _10608_ (
    .A1(_00150_),
    .A2(_00151_),
    .B1(addr_i_3_),
    .Y(_00152_)
  );
  sg13g2_a22oi_1 _10609_ (
    .A1(_00146_),
    .A2(_00149_),
    .B1(_00152_),
    .B2(_07403_),
    .Y(_00153_)
  );
  sg13g2_buf_1 _10610_ (
    .A(_01066_),
    .X(_00155_)
  );
  sg13g2_buf_1 _10611_ (
    .A(_08111_),
    .X(_00156_)
  );
  sg13g2_buf_1 _10612_ (
    .A(_00319_),
    .X(_00157_)
  );
  sg13g2_buf_1 _10613_ (
    .A(_04937_),
    .X(_00158_)
  );
  sg13g2_buf_1 _10614_ (
    .A(_00158_),
    .X(_00159_)
  );
  sg13g2_a22oi_1 _10615_ (
    .A1(_00155_),
    .A2(_00156_),
    .B1(_00157_),
    .B2(_00159_),
    .Y(_00160_)
  );
  sg13g2_nand2b_1 _10616_ (
    .A_N(_00160_),
    .B(addr_i_5_),
    .Y(_00161_)
  );
  sg13g2_a21oi_1 _10617_ (
    .A1(_00153_),
    .A2(_00161_),
    .B1(_03073_),
    .Y(_00162_)
  );
  sg13g2_o21ai_1 _10618_ (
    .A1(_03238_),
    .A2(_00144_),
    .B1(_00162_),
    .Y(_00163_)
  );
  sg13g2_a22oi_1 _10619_ (
    .A1(_00114_),
    .A2(_00130_),
    .B1(_00135_),
    .B2(_00163_),
    .Y(_00164_)
  );
  sg13g2_a22oi_1 _10620_ (
    .A1(_09490_),
    .A2(_00045_),
    .B1(_00111_),
    .B2(_00164_),
    .Y(_00166_)
  );
  sg13g2_nor2_1 _10621_ (
    .A(addr_i_11_),
    .B(_00166_),
    .Y(_00167_)
  );
  sg13g2_buf_1 _10622_ (
    .A(_02623_),
    .X(_00168_)
  );
  sg13g2_buf_1 _10623_ (
    .A(_00168_),
    .X(_00169_)
  );
  sg13g2_nor2_1 _10624_ (
    .A(addr_i_4_),
    .B(addr_i_8_),
    .Y(_00170_)
  );
  sg13g2_nand2_1 _10625_ (
    .A(_00170_),
    .B(_07911_),
    .Y(_00171_)
  );
  sg13g2_buf_1 _10626_ (
    .A(_06717_),
    .X(_00172_)
  );
  sg13g2_nand2_1 _10627_ (
    .A(_03765_),
    .B(_08564_),
    .Y(_00173_)
  );
  sg13g2_o21ai_1 _10628_ (
    .A1(addr_i_3_),
    .A2(_00173_),
    .B1(_05490_),
    .Y(_00174_)
  );
  sg13g2_and3_1 _10629_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .C(addr_i_5_),
    .X(_00175_)
  );
  sg13g2_buf_1 _10630_ (
    .A(_00175_),
    .X(_00177_)
  );
  sg13g2_o21ai_1 _10631_ (
    .A1(_06806_),
    .A2(_00177_),
    .B1(addr_i_3_),
    .Y(_00178_)
  );
  sg13g2_a22oi_1 _10632_ (
    .A1(_00022_),
    .A2(_05535_),
    .B1(_01285_),
    .B2(_09094_),
    .Y(_00179_)
  );
  sg13g2_nand2_1 _10633_ (
    .A(_00178_),
    .B(_00179_),
    .Y(_00180_)
  );
  sg13g2_a21oi_1 _10634_ (
    .A1(_00172_),
    .A2(_00174_),
    .B1(_00180_),
    .Y(_00181_)
  );
  sg13g2_a22oi_1 _10635_ (
    .A1(_00169_),
    .A2(_00171_),
    .B1(_00181_),
    .B2(addr_i_9_),
    .Y(_00182_)
  );
  sg13g2_buf_1 _10636_ (
    .A(_09501_),
    .X(_00183_)
  );
  sg13g2_o21ai_1 _10637_ (
    .A1(addr_i_2_),
    .A2(addr_i_5_),
    .B1(addr_i_6_),
    .Y(_00184_)
  );
  sg13g2_buf_1 _10638_ (
    .A(_08796_),
    .X(_00185_)
  );
  sg13g2_nand2_1 _10639_ (
    .A(_03270_),
    .B(_08597_),
    .Y(_00186_)
  );
  sg13g2_a21oi_1 _10640_ (
    .A1(_00185_),
    .A2(_00186_),
    .B1(addr_i_4_),
    .Y(_00188_)
  );
  sg13g2_a22oi_1 _10641_ (
    .A1(_00183_),
    .A2(_00184_),
    .B1(_00188_),
    .B2(addr_i_3_),
    .Y(_00189_)
  );
  sg13g2_buf_1 _10642_ (
    .A(_08785_),
    .X(_00190_)
  );
  sg13g2_buf_1 _10643_ (
    .A(_00190_),
    .X(_00191_)
  );
  sg13g2_buf_1 _10644_ (
    .A(_03523_),
    .X(_00192_)
  );
  sg13g2_nor3_1 _10645_ (
    .A(_00191_),
    .B(_06950_),
    .C(_00192_),
    .Y(_00193_)
  );
  sg13g2_xnor2_1 _10646_ (
    .A(addr_i_4_),
    .B(addr_i_7_),
    .Y(_00194_)
  );
  sg13g2_nand2_1 _10647_ (
    .A(_07558_),
    .B(_09478_),
    .Y(_00195_)
  );
  sg13g2_a22oi_1 _10648_ (
    .A1(_00194_),
    .A2(_00195_),
    .B1(addr_i_8_),
    .B2(_00169_),
    .Y(_00196_)
  );
  sg13g2_o21ai_1 _10649_ (
    .A1(_00189_),
    .A2(_00193_),
    .B1(_00196_),
    .Y(_00197_)
  );
  sg13g2_buf_1 _10650_ (
    .A(_03435_),
    .X(_00199_)
  );
  sg13g2_buf_1 _10651_ (
    .A(_00199_),
    .X(_00200_)
  );
  sg13g2_nor2_1 _10652_ (
    .A(_00200_),
    .B(_01011_),
    .Y(_00201_)
  );
  sg13g2_a21oi_1 _10653_ (
    .A1(addr_i_6_),
    .A2(_03238_),
    .B1(_00201_),
    .Y(_00202_)
  );
  sg13g2_a221oi_1 _10654_ (
    .A1(_00182_),
    .A2(_00197_),
    .B1(_00202_),
    .B2(addr_i_9_),
    .C1(addr_i_10_),
    .Y(_00203_)
  );
  sg13g2_a21oi_1 _10655_ (
    .A1(_06485_),
    .A2(_07713_),
    .B1(addr_i_3_),
    .Y(_00204_)
  );
  sg13g2_nor2_1 _10656_ (
    .A(addr_i_4_),
    .B(_06485_),
    .Y(_00205_)
  );
  sg13g2_buf_1 _10657_ (
    .A(_00205_),
    .X(_00206_)
  );
  sg13g2_o21ai_1 _10658_ (
    .A1(_00204_),
    .A2(_00206_),
    .B1(addr_i_2_),
    .Y(_00207_)
  );
  sg13g2_nor2b_1 _10659_ (
    .A(addr_i_2_),
    .B_N(addr_i_3_),
    .Y(_00208_)
  );
  sg13g2_buf_1 _10660_ (
    .A(_00208_),
    .X(_00210_)
  );
  sg13g2_nand2_1 _10661_ (
    .A(_00539_),
    .B(_00210_),
    .Y(_00211_)
  );
  sg13g2_nand3_1 _10662_ (
    .A(addr_i_7_),
    .B(_00207_),
    .C(_00211_),
    .Y(_00212_)
  );
  sg13g2_nand2_1 _10663_ (
    .A(_00374_),
    .B(_01537_),
    .Y(_00213_)
  );
  sg13g2_buf_1 _10664_ (
    .A(_00213_),
    .X(_00214_)
  );
  sg13g2_nor2_1 _10665_ (
    .A(_03731_),
    .B(_00214_),
    .Y(_00215_)
  );
  sg13g2_nand3_1 _10666_ (
    .A(_00069_),
    .B(_00212_),
    .C(_00215_),
    .Y(_00216_)
  );
  sg13g2_nand2_1 _10667_ (
    .A(addr_i_11_),
    .B(_00216_),
    .Y(_00217_)
  );
  sg13g2_o21ai_1 _10668_ (
    .A1(_00203_),
    .A2(_00217_),
    .B1(addr_i_12_),
    .Y(_00218_)
  );
  sg13g2_a21oi_1 _10669_ (
    .A1(addr_i_5_),
    .A2(_00890_),
    .B1(_04849_),
    .Y(_00219_)
  );
  sg13g2_nor2_1 _10670_ (
    .A(_00191_),
    .B(_00219_),
    .Y(_00221_)
  );
  sg13g2_nor3_1 _10671_ (
    .A(_04683_),
    .B(_02963_),
    .C(_00221_),
    .Y(_00222_)
  );
  sg13g2_buf_1 _10672_ (
    .A(_04119_),
    .X(_00223_)
  );
  sg13g2_nand2_1 _10673_ (
    .A(_09038_),
    .B(_07956_),
    .Y(_00224_)
  );
  sg13g2_o21ai_1 _10674_ (
    .A1(_00223_),
    .A2(_07889_),
    .B1(_00224_),
    .Y(_00225_)
  );
  sg13g2_nor2_1 _10675_ (
    .A(_07933_),
    .B(_00462_),
    .Y(_00226_)
  );
  sg13g2_buf_1 _10676_ (
    .A(_00226_),
    .X(_00227_)
  );
  sg13g2_nand2_1 _10677_ (
    .A(_03446_),
    .B(_04528_),
    .Y(_00228_)
  );
  sg13g2_a21oi_1 _10678_ (
    .A1(_02810_),
    .A2(_00228_),
    .B1(addr_i_3_),
    .Y(_00229_)
  );
  sg13g2_buf_1 _10679_ (
    .A(_02569_),
    .X(_00230_)
  );
  sg13g2_a22oi_1 _10680_ (
    .A1(addr_i_3_),
    .A2(_00227_),
    .B1(_00229_),
    .B2(_00230_),
    .Y(_00232_)
  );
  sg13g2_a22oi_1 _10681_ (
    .A1(_09138_),
    .A2(_00225_),
    .B1(_00232_),
    .B2(addr_i_8_),
    .Y(_00233_)
  );
  sg13g2_nor2_1 _10682_ (
    .A(addr_i_7_),
    .B(_05734_),
    .Y(_00234_)
  );
  sg13g2_o21ai_1 _10683_ (
    .A1(_00110_),
    .A2(_08144_),
    .B1(addr_i_3_),
    .Y(_00235_)
  );
  sg13g2_inv_1 _10684_ (
    .A(_00235_),
    .Y(_00236_)
  );
  sg13g2_o21ai_1 _10685_ (
    .A1(_00234_),
    .A2(_00236_),
    .B1(addr_i_5_),
    .Y(_00237_)
  );
  sg13g2_buf_1 _10686_ (
    .A(_00208_),
    .X(_00238_)
  );
  sg13g2_buf_1 _10687_ (
    .A(_00238_),
    .X(_00239_)
  );
  sg13g2_o21ai_1 _10688_ (
    .A1(_06740_),
    .A2(_00239_),
    .B1(_07889_),
    .Y(_00240_)
  );
  sg13g2_nand3_1 _10689_ (
    .A(_07038_),
    .B(_00237_),
    .C(_00240_),
    .Y(_00241_)
  );
  sg13g2_buf_1 _10690_ (
    .A(_00385_),
    .X(_00243_)
  );
  sg13g2_buf_1 _10691_ (
    .A(_03194_),
    .X(_00244_)
  );
  sg13g2_nand2b_1 _10692_ (
    .A_N(addr_i_2_),
    .B(addr_i_7_),
    .Y(_00245_)
  );
  sg13g2_buf_1 _10693_ (
    .A(_00245_),
    .X(_00246_)
  );
  sg13g2_nor2_1 _10694_ (
    .A(addr_i_4_),
    .B(_00246_),
    .Y(_00247_)
  );
  sg13g2_o21ai_1 _10695_ (
    .A1(_00244_),
    .A2(_00247_),
    .B1(addr_i_3_),
    .Y(_00248_)
  );
  sg13g2_nand2_1 _10696_ (
    .A(_00044_),
    .B(_06729_),
    .Y(_00249_)
  );
  sg13g2_nand2_1 _10697_ (
    .A(addr_i_4_),
    .B(_00154_),
    .Y(_00250_)
  );
  sg13g2_a21oi_1 _10698_ (
    .A1(_00249_),
    .A2(_00250_),
    .B1(addr_i_3_),
    .Y(_00251_)
  );
  sg13g2_buf_1 _10699_ (
    .A(_07956_),
    .X(_00252_)
  );
  sg13g2_nor2_1 _10700_ (
    .A(addr_i_7_),
    .B(_00252_),
    .Y(_00254_)
  );
  sg13g2_nor2_1 _10701_ (
    .A(addr_i_5_),
    .B(_00254_),
    .Y(_00255_)
  );
  sg13g2_nor4_1 _10702_ (
    .A(addr_i_6_),
    .B(_00017_),
    .C(_00251_),
    .D(_00255_),
    .Y(_00256_)
  );
  sg13g2_nor2_1 _10703_ (
    .A(addr_i_2_),
    .B(_02272_),
    .Y(_00257_)
  );
  sg13g2_buf_1 _10704_ (
    .A(_08111_),
    .X(_00258_)
  );
  sg13g2_o21ai_1 _10705_ (
    .A1(_09061_),
    .A2(_00257_),
    .B1(_00258_),
    .Y(_00259_)
  );
  sg13g2_buf_1 _10706_ (
    .A(_07491_),
    .X(_00260_)
  );
  sg13g2_buf_1 _10707_ (
    .A(_00260_),
    .X(_00261_)
  );
  sg13g2_buf_1 _10708_ (
    .A(_04284_),
    .X(_00262_)
  );
  sg13g2_o21ai_1 _10709_ (
    .A1(_00261_),
    .A2(_07503_),
    .B1(_00262_),
    .Y(_00263_)
  );
  sg13g2_a21oi_1 _10710_ (
    .A1(_00259_),
    .A2(_00263_),
    .B1(addr_i_5_),
    .Y(_00265_)
  );
  sg13g2_nor2_1 _10711_ (
    .A(_07049_),
    .B(_08863_),
    .Y(_00266_)
  );
  sg13g2_nand3b_1 _10712_ (
    .A_N(_00266_),
    .B(_00168_),
    .C(_09476_),
    .Y(_00267_)
  );
  sg13g2_buf_1 _10713_ (
    .A(_08166_),
    .X(_00268_)
  );
  sg13g2_buf_1 _10714_ (
    .A(_08885_),
    .X(_00269_)
  );
  sg13g2_nor3_1 _10715_ (
    .A(addr_i_3_),
    .B(_00269_),
    .C(_08144_),
    .Y(_00270_)
  );
  sg13g2_o21ai_1 _10716_ (
    .A1(_00268_),
    .A2(_00270_),
    .B1(_05247_),
    .Y(_00271_)
  );
  sg13g2_nand3_1 _10717_ (
    .A(addr_i_8_),
    .B(_00267_),
    .C(_00271_),
    .Y(_00272_)
  );
  sg13g2_a22oi_1 _10718_ (
    .A1(_00248_),
    .A2(_00256_),
    .B1(_00265_),
    .B2(_00272_),
    .Y(_00273_)
  );
  sg13g2_a22oi_1 _10719_ (
    .A1(_00233_),
    .A2(_00241_),
    .B1(_00243_),
    .B2(_00273_),
    .Y(_00274_)
  );
  sg13g2_buf_1 _10720_ (
    .A(_04650_),
    .X(_00276_)
  );
  sg13g2_buf_1 _10721_ (
    .A(_00276_),
    .X(_00277_)
  );
  sg13g2_nor2_1 _10722_ (
    .A(addr_i_3_),
    .B(_00462_),
    .Y(_00278_)
  );
  sg13g2_buf_1 _10723_ (
    .A(_00278_),
    .X(_00279_)
  );
  sg13g2_nor2_1 _10724_ (
    .A(_01757_),
    .B(_08941_),
    .Y(_00280_)
  );
  sg13g2_or2_1 _10725_ (
    .A(_00279_),
    .B(_00280_),
    .X(_00281_)
  );
  sg13g2_nor2_1 _10726_ (
    .A(_03270_),
    .B(_00835_),
    .Y(_00282_)
  );
  sg13g2_nand2_1 _10727_ (
    .A(_00258_),
    .B(_00282_),
    .Y(_00283_)
  );
  sg13g2_buf_1 _10728_ (
    .A(_03490_),
    .X(_00284_)
  );
  sg13g2_a21oi_1 _10729_ (
    .A1(_04715_),
    .A2(_00284_),
    .B1(addr_i_3_),
    .Y(_00285_)
  );
  sg13g2_nand3_1 _10730_ (
    .A(addr_i_3_),
    .B(addr_i_2_),
    .C(addr_i_5_),
    .Y(_00287_)
  );
  sg13g2_a21oi_1 _10731_ (
    .A1(_04162_),
    .A2(_00287_),
    .B1(addr_i_6_),
    .Y(_00288_)
  );
  sg13g2_o21ai_1 _10732_ (
    .A1(_00285_),
    .A2(_00288_),
    .B1(_09271_),
    .Y(_00289_)
  );
  sg13g2_buf_1 _10733_ (
    .A(_01494_),
    .X(_00290_)
  );
  sg13g2_a21oi_1 _10734_ (
    .A1(_00283_),
    .A2(_00289_),
    .B1(_00290_),
    .Y(_00291_)
  );
  sg13g2_buf_1 _10735_ (
    .A(_07061_),
    .X(_00292_)
  );
  sg13g2_buf_1 _10736_ (
    .A(_03446_),
    .X(_00293_)
  );
  sg13g2_buf_1 _10737_ (
    .A(_06729_),
    .X(_00294_)
  );
  sg13g2_nor3_1 _10738_ (
    .A(_04041_),
    .B(_00293_),
    .C(_00294_),
    .Y(_00295_)
  );
  sg13g2_o21ai_1 _10739_ (
    .A1(_00292_),
    .A2(_00295_),
    .B1(addr_i_4_),
    .Y(_00296_)
  );
  sg13g2_buf_1 _10740_ (
    .A(_05524_),
    .X(_00298_)
  );
  sg13g2_o21ai_1 _10741_ (
    .A1(addr_i_5_),
    .A2(_04173_),
    .B1(_04793_),
    .Y(_00299_)
  );
  sg13g2_a21oi_1 _10742_ (
    .A1(_00298_),
    .A2(_00299_),
    .B1(_00060_),
    .Y(_00300_)
  );
  sg13g2_buf_1 _10743_ (
    .A(_03643_),
    .X(_00301_)
  );
  sg13g2_nand2_1 _10744_ (
    .A(addr_i_7_),
    .B(_00024_),
    .Y(_00302_)
  );
  sg13g2_nor2b_1 _10745_ (
    .A(addr_i_6_),
    .B_N(addr_i_4_),
    .Y(_00303_)
  );
  sg13g2_buf_1 _10746_ (
    .A(_00303_),
    .X(_00304_)
  );
  sg13g2_buf_1 _10747_ (
    .A(_00304_),
    .X(_00305_)
  );
  sg13g2_a221oi_1 _10748_ (
    .A1(_00298_),
    .A2(_00301_),
    .B1(_00302_),
    .B2(_00305_),
    .C1(addr_i_3_),
    .Y(_00306_)
  );
  sg13g2_a22oi_1 _10749_ (
    .A1(_00296_),
    .A2(_00300_),
    .B1(_00306_),
    .B2(addr_i_8_),
    .Y(_00307_)
  );
  sg13g2_a22oi_1 _10750_ (
    .A1(_00277_),
    .A2(_00281_),
    .B1(_00291_),
    .B2(_00307_),
    .Y(_00309_)
  );
  sg13g2_nor2_1 _10751_ (
    .A(addr_i_9_),
    .B(_00309_),
    .Y(_00310_)
  );
  sg13g2_nor4_1 _10752_ (
    .A(addr_i_10_),
    .B(_00222_),
    .C(_00274_),
    .D(_00310_),
    .Y(_00311_)
  );
  sg13g2_nor2_1 _10753_ (
    .A(addr_i_12_),
    .B(addr_i_11_),
    .Y(_00312_)
  );
  sg13g2_nor2b_1 _10754_ (
    .A(_00311_),
    .B_N(_00312_),
    .Y(_00313_)
  );
  sg13g2_nand2_1 _10755_ (
    .A(_05346_),
    .B(_02645_),
    .Y(_00314_)
  );
  sg13g2_buf_1 _10756_ (
    .A(_08464_),
    .X(_00315_)
  );
  sg13g2_buf_1 _10757_ (
    .A(_02547_),
    .X(_00316_)
  );
  sg13g2_buf_1 _10758_ (
    .A(_00316_),
    .X(_00317_)
  );
  sg13g2_a22oi_1 _10759_ (
    .A1(addr_i_4_),
    .A2(_00315_),
    .B1(_00317_),
    .B2(_00015_),
    .Y(_00318_)
  );
  sg13g2_nand2_1 _10760_ (
    .A(addr_i_2_),
    .B(_01197_),
    .Y(_00320_)
  );
  sg13g2_nand2_1 _10761_ (
    .A(_04373_),
    .B(_00320_),
    .Y(_00321_)
  );
  sg13g2_buf_1 _10762_ (
    .A(_04218_),
    .X(_00322_)
  );
  sg13g2_o21ai_1 _10763_ (
    .A1(addr_i_5_),
    .A2(_00322_),
    .B1(addr_i_4_),
    .Y(_00323_)
  );
  sg13g2_buf_1 _10764_ (
    .A(_00021_),
    .X(_00324_)
  );
  sg13g2_a21oi_1 _10765_ (
    .A1(_00321_),
    .A2(_00323_),
    .B1(_00324_),
    .Y(_00325_)
  );
  sg13g2_a22oi_1 _10766_ (
    .A1(_00314_),
    .A2(_00318_),
    .B1(_00325_),
    .B2(addr_i_8_),
    .Y(_00326_)
  );
  sg13g2_buf_1 _10767_ (
    .A(_07469_),
    .X(_00327_)
  );
  sg13g2_nand2_1 _10768_ (
    .A(_00117_),
    .B(_00327_),
    .Y(_00328_)
  );
  sg13g2_nor2_1 _10769_ (
    .A(addr_i_2_),
    .B(_04860_),
    .Y(_00329_)
  );
  sg13g2_o21ai_1 _10770_ (
    .A1(addr_i_3_),
    .A2(_00329_),
    .B1(_00155_),
    .Y(_00331_)
  );
  sg13g2_a22oi_1 _10771_ (
    .A1(addr_i_3_),
    .A2(_00328_),
    .B1(_00331_),
    .B2(_00659_),
    .Y(_00332_)
  );
  sg13g2_nand2_1 _10772_ (
    .A(addr_i_3_),
    .B(addr_i_6_),
    .Y(_00333_)
  );
  sg13g2_nor2_1 _10773_ (
    .A(addr_i_5_),
    .B(_00333_),
    .Y(_00334_)
  );
  sg13g2_a21oi_1 _10774_ (
    .A1(addr_i_5_),
    .A2(_03743_),
    .B1(addr_i_2_),
    .Y(_00335_)
  );
  sg13g2_nor3_1 _10775_ (
    .A(addr_i_4_),
    .B(_00334_),
    .C(_00335_),
    .Y(_00336_)
  );
  sg13g2_o21ai_1 _10776_ (
    .A1(_00332_),
    .A2(_00336_),
    .B1(addr_i_7_),
    .Y(_00337_)
  );
  sg13g2_nor2_1 _10777_ (
    .A(addr_i_4_),
    .B(_00038_),
    .Y(_00338_)
  );
  sg13g2_buf_1 _10778_ (
    .A(_01834_),
    .X(_00339_)
  );
  sg13g2_nand2_1 _10779_ (
    .A(_00190_),
    .B(_00339_),
    .Y(_00340_)
  );
  sg13g2_buf_1 _10780_ (
    .A(_00033_),
    .X(_00342_)
  );
  sg13g2_buf_1 _10781_ (
    .A(_00342_),
    .X(_00343_)
  );
  sg13g2_o21ai_1 _10782_ (
    .A1(_00343_),
    .A2(_08653_),
    .B1(addr_i_3_),
    .Y(_00344_)
  );
  sg13g2_o21ai_1 _10783_ (
    .A1(_00338_),
    .A2(_00340_),
    .B1(_00344_),
    .Y(_00345_)
  );
  sg13g2_nor2_1 _10784_ (
    .A(addr_i_3_),
    .B(_01625_),
    .Y(_00346_)
  );
  sg13g2_buf_1 _10785_ (
    .A(_05700_),
    .X(_00347_)
  );
  sg13g2_nor2_1 _10786_ (
    .A(_00347_),
    .B(_06032_),
    .Y(_00348_)
  );
  sg13g2_o21ai_1 _10787_ (
    .A1(_00346_),
    .A2(_00348_),
    .B1(_05600_),
    .Y(_00349_)
  );
  sg13g2_nand2_1 _10788_ (
    .A(addr_i_8_),
    .B(_00349_),
    .Y(_00350_)
  );
  sg13g2_buf_1 _10789_ (
    .A(_05811_),
    .X(_00351_)
  );
  sg13g2_buf_1 _10790_ (
    .A(_09415_),
    .X(_00353_)
  );
  sg13g2_buf_1 _10791_ (
    .A(_00044_),
    .X(_00354_)
  );
  sg13g2_nand2_1 _10792_ (
    .A(_00354_),
    .B(_00184_),
    .Y(_00355_)
  );
  sg13g2_a21oi_1 _10793_ (
    .A1(_00353_),
    .A2(_00355_),
    .B1(addr_i_3_),
    .Y(_00356_)
  );
  sg13g2_nand3b_1 _10794_ (
    .A_N(addr_i_3_),
    .B(addr_i_2_),
    .C(addr_i_6_),
    .Y(_00357_)
  );
  sg13g2_buf_1 _10795_ (
    .A(_00357_),
    .X(_00358_)
  );
  sg13g2_nand3_1 _10796_ (
    .A(addr_i_3_),
    .B(addr_i_5_),
    .C(_08774_),
    .Y(_00359_)
  );
  sg13g2_buf_1 _10797_ (
    .A(_00354_),
    .X(_00360_)
  );
  sg13g2_a21oi_1 _10798_ (
    .A1(_00358_),
    .A2(_00359_),
    .B1(_00360_),
    .Y(_00361_)
  );
  sg13g2_nor4_1 _10799_ (
    .A(_00351_),
    .B(_03501_),
    .C(_00356_),
    .D(_00361_),
    .Y(_00362_)
  );
  sg13g2_a22oi_1 _10800_ (
    .A1(_09474_),
    .A2(_00345_),
    .B1(_00350_),
    .B2(_00362_),
    .Y(_00364_)
  );
  sg13g2_a21oi_1 _10801_ (
    .A1(_00326_),
    .A2(_00337_),
    .B1(_00364_),
    .Y(_00365_)
  );
  sg13g2_nand2_1 _10802_ (
    .A(addr_i_9_),
    .B(_00365_),
    .Y(_00366_)
  );
  sg13g2_buf_1 _10803_ (
    .A(_05888_),
    .X(_00367_)
  );
  sg13g2_nand2_1 _10804_ (
    .A(addr_i_4_),
    .B(_00000_),
    .Y(_00368_)
  );
  sg13g2_a21oi_1 _10805_ (
    .A1(_01757_),
    .A2(_00368_),
    .B1(_08156_),
    .Y(_00369_)
  );
  sg13g2_nand2_1 _10806_ (
    .A(_00033_),
    .B(_00539_),
    .Y(_00370_)
  );
  sg13g2_buf_1 _10807_ (
    .A(_00370_),
    .X(_00371_)
  );
  sg13g2_a21oi_1 _10808_ (
    .A1(_00371_),
    .A2(_02634_),
    .B1(addr_i_3_),
    .Y(_00372_)
  );
  sg13g2_o21ai_1 _10809_ (
    .A1(_00369_),
    .A2(_00372_),
    .B1(_06619_),
    .Y(_00373_)
  );
  sg13g2_buf_1 _10810_ (
    .A(_03665_),
    .X(_00375_)
  );
  sg13g2_buf_1 _10811_ (
    .A(_00303_),
    .X(_00376_)
  );
  sg13g2_buf_1 _10812_ (
    .A(_05169_),
    .X(_00377_)
  );
  sg13g2_o21ai_1 _10813_ (
    .A1(_00375_),
    .A2(_00376_),
    .B1(_00377_),
    .Y(_00378_)
  );
  sg13g2_a21oi_1 _10814_ (
    .A1(_00373_),
    .A2(_00378_),
    .B1(_03292_),
    .Y(_00379_)
  );
  sg13g2_buf_1 _10815_ (
    .A(_03952_),
    .X(_00380_)
  );
  sg13g2_buf_1 _10816_ (
    .A(_00380_),
    .X(_00381_)
  );
  sg13g2_nand3_1 _10817_ (
    .A(addr_i_7_),
    .B(_00381_),
    .C(_06873_),
    .Y(_00382_)
  );
  sg13g2_nor2b_1 _10818_ (
    .A(addr_i_4_),
    .B_N(addr_i_7_),
    .Y(_00383_)
  );
  sg13g2_buf_1 _10819_ (
    .A(_00383_),
    .X(_00384_)
  );
  sg13g2_buf_1 _10820_ (
    .A(_00384_),
    .X(_00386_)
  );
  sg13g2_o21ai_1 _10821_ (
    .A1(_00386_),
    .A2(_05568_),
    .B1(addr_i_3_),
    .Y(_00387_)
  );
  sg13g2_buf_1 _10822_ (
    .A(_02777_),
    .X(_00388_)
  );
  sg13g2_a21oi_1 _10823_ (
    .A1(_00382_),
    .A2(_00387_),
    .B1(_00388_),
    .Y(_00389_)
  );
  sg13g2_buf_1 _10824_ (
    .A(_02569_),
    .X(_00390_)
  );
  sg13g2_buf_1 _10825_ (
    .A(_02250_),
    .X(_00391_)
  );
  sg13g2_a21oi_1 _10826_ (
    .A1(_00390_),
    .A2(_03358_),
    .B1(_00391_),
    .Y(_00392_)
  );
  sg13g2_nor4_1 _10827_ (
    .A(_00367_),
    .B(_00379_),
    .C(_00389_),
    .D(_00392_),
    .Y(_00393_)
  );
  sg13g2_nand2_1 _10828_ (
    .A(_09459_),
    .B(_07503_),
    .Y(_00394_)
  );
  sg13g2_nor2_1 _10829_ (
    .A(_03062_),
    .B(_00394_),
    .Y(_00395_)
  );
  sg13g2_buf_1 _10830_ (
    .A(_02700_),
    .X(_00397_)
  );
  sg13g2_o21ai_1 _10831_ (
    .A1(_00393_),
    .A2(_00395_),
    .B1(_00397_),
    .Y(_00398_)
  );
  sg13g2_nor2_1 _10832_ (
    .A(_08564_),
    .B(_00198_),
    .Y(_00399_)
  );
  sg13g2_buf_1 _10833_ (
    .A(_07237_),
    .X(_00400_)
  );
  sg13g2_buf_1 _10834_ (
    .A(_00400_),
    .X(_00401_)
  );
  sg13g2_buf_1 _10835_ (
    .A(_09486_),
    .X(_00402_)
  );
  sg13g2_buf_1 _10836_ (
    .A(_08930_),
    .X(_00403_)
  );
  sg13g2_nand2_1 _10837_ (
    .A(_04550_),
    .B(_00066_),
    .Y(_00404_)
  );
  sg13g2_buf_1 _10838_ (
    .A(_00404_),
    .X(_00405_)
  );
  sg13g2_buf_1 _10839_ (
    .A(_00078_),
    .X(_00406_)
  );
  sg13g2_buf_1 _10840_ (
    .A(_00406_),
    .X(_00408_)
  );
  sg13g2_buf_1 _10841_ (
    .A(_00408_),
    .X(_00409_)
  );
  sg13g2_a21oi_1 _10842_ (
    .A1(_00403_),
    .A2(_00405_),
    .B1(_00409_),
    .Y(_00410_)
  );
  sg13g2_a22oi_1 _10843_ (
    .A1(_00401_),
    .A2(_00402_),
    .B1(_07215_),
    .B2(_00410_),
    .Y(_00411_)
  );
  sg13g2_nor2_1 _10844_ (
    .A(addr_i_6_),
    .B(_09493_),
    .Y(_00412_)
  );
  sg13g2_buf_1 _10845_ (
    .A(_03490_),
    .X(_00413_)
  );
  sg13g2_buf_1 _10846_ (
    .A(_00413_),
    .X(_00414_)
  );
  sg13g2_nor2_1 _10847_ (
    .A(addr_i_4_),
    .B(_00495_),
    .Y(_00415_)
  );
  sg13g2_nor2_1 _10848_ (
    .A(_01581_),
    .B(_00406_),
    .Y(_00416_)
  );
  sg13g2_nor2_1 _10849_ (
    .A(_00415_),
    .B(_00416_),
    .Y(_00417_)
  );
  sg13g2_a21oi_1 _10850_ (
    .A1(_00414_),
    .A2(_00417_),
    .B1(addr_i_7_),
    .Y(_00419_)
  );
  sg13g2_a22oi_1 _10851_ (
    .A1(_06740_),
    .A2(_00412_),
    .B1(_00419_),
    .B2(addr_i_3_),
    .Y(_00420_)
  );
  sg13g2_a21oi_1 _10852_ (
    .A1(addr_i_3_),
    .A2(_00411_),
    .B1(_00420_),
    .Y(_00421_)
  );
  sg13g2_nor2_1 _10853_ (
    .A(addr_i_9_),
    .B(addr_i_8_),
    .Y(_00422_)
  );
  sg13g2_buf_1 _10854_ (
    .A(_00422_),
    .X(_00423_)
  );
  sg13g2_o21ai_1 _10855_ (
    .A1(_00399_),
    .A2(_00421_),
    .B1(_00423_),
    .Y(_00424_)
  );
  sg13g2_nand4_1 _10856_ (
    .A(addr_i_10_),
    .B(_00366_),
    .C(_00398_),
    .D(_00424_),
    .Y(_00425_)
  );
  sg13g2_nor2_1 _10857_ (
    .A(_06496_),
    .B(_08885_),
    .Y(_00426_)
  );
  sg13g2_nand2_1 _10858_ (
    .A(_09050_),
    .B(_00252_),
    .Y(_00427_)
  );
  sg13g2_buf_1 _10859_ (
    .A(_02623_),
    .X(_00428_)
  );
  sg13g2_nand2_1 _10860_ (
    .A(_00120_),
    .B(_03380_),
    .Y(_00430_)
  );
  sg13g2_nand3_1 _10861_ (
    .A(_00428_),
    .B(_01208_),
    .C(_00430_),
    .Y(_00431_)
  );
  sg13g2_nand3_1 _10862_ (
    .A(addr_i_8_),
    .B(_00427_),
    .C(_00431_),
    .Y(_00432_)
  );
  sg13g2_nand2_1 _10863_ (
    .A(addr_i_2_),
    .B(_04173_),
    .Y(_00433_)
  );
  sg13g2_buf_1 _10864_ (
    .A(_00433_),
    .X(_00434_)
  );
  sg13g2_buf_1 _10865_ (
    .A(_02272_),
    .X(_00435_)
  );
  sg13g2_nor2_1 _10866_ (
    .A(_00435_),
    .B(_05457_),
    .Y(_00436_)
  );
  sg13g2_o21ai_1 _10867_ (
    .A1(_09061_),
    .A2(_00436_),
    .B1(addr_i_3_),
    .Y(_00437_)
  );
  sg13g2_a21oi_1 _10868_ (
    .A1(_00434_),
    .A2(_00437_),
    .B1(addr_i_5_),
    .Y(_00438_)
  );
  sg13g2_a22oi_1 _10869_ (
    .A1(_00183_),
    .A2(_00426_),
    .B1(_00432_),
    .B2(_00438_),
    .Y(_00439_)
  );
  sg13g2_buf_1 _10870_ (
    .A(_04075_),
    .X(_00441_)
  );
  sg13g2_buf_1 _10871_ (
    .A(_02645_),
    .X(_00442_)
  );
  sg13g2_nand2_1 _10872_ (
    .A(_00441_),
    .B(_00442_),
    .Y(_00443_)
  );
  sg13g2_a21o_1 _10873_ (
    .A1(_04639_),
    .A2(_00443_),
    .B1(_00230_),
    .X(_00444_)
  );
  sg13g2_buf_1 _10874_ (
    .A(_00199_),
    .X(_00445_)
  );
  sg13g2_o21ai_1 _10875_ (
    .A1(addr_i_2_),
    .A2(_00383_),
    .B1(_09393_),
    .Y(_00446_)
  );
  sg13g2_xnor2_1 _10876_ (
    .A(addr_i_2_),
    .B(addr_i_6_),
    .Y(_00447_)
  );
  sg13g2_buf_1 _10877_ (
    .A(_00447_),
    .X(_00448_)
  );
  sg13g2_nor2_1 _10878_ (
    .A(_02602_),
    .B(_00448_),
    .Y(_00449_)
  );
  sg13g2_a21oi_1 _10879_ (
    .A1(_00445_),
    .A2(_00446_),
    .B1(_00449_),
    .Y(_00450_)
  );
  sg13g2_or2_1 _10880_ (
    .A(addr_i_3_),
    .B(_00450_),
    .X(_00452_)
  );
  sg13g2_nand2_1 _10881_ (
    .A(_03908_),
    .B(_00154_),
    .Y(_00453_)
  );
  sg13g2_buf_1 _10882_ (
    .A(_05722_),
    .X(_00454_)
  );
  sg13g2_o21ai_1 _10883_ (
    .A1(_00454_),
    .A2(_00158_),
    .B1(addr_i_4_),
    .Y(_00455_)
  );
  sg13g2_nand3_1 _10884_ (
    .A(_00434_),
    .B(_00453_),
    .C(_00455_),
    .Y(_00456_)
  );
  sg13g2_a22oi_1 _10885_ (
    .A1(addr_i_3_),
    .A2(_00456_),
    .B1(_05600_),
    .B2(_04439_),
    .Y(_00457_)
  );
  sg13g2_nand2_1 _10886_ (
    .A(_04151_),
    .B(_08343_),
    .Y(_00458_)
  );
  sg13g2_and4_1 _10887_ (
    .A(_05600_),
    .B(_01921_),
    .C(_09476_),
    .D(_00458_),
    .X(_00459_)
  );
  sg13g2_a22oi_1 _10888_ (
    .A1(_00452_),
    .A2(_00457_),
    .B1(addr_i_8_),
    .B2(_00459_),
    .Y(_00460_)
  );
  sg13g2_a21oi_1 _10889_ (
    .A1(_00439_),
    .A2(_00444_),
    .B1(_00460_),
    .Y(_00461_)
  );
  sg13g2_buf_1 _10890_ (
    .A(_05845_),
    .X(_00463_)
  );
  sg13g2_o21ai_1 _10891_ (
    .A1(addr_i_4_),
    .A2(_05335_),
    .B1(_00019_),
    .Y(_00464_)
  );
  sg13g2_and2_1 _10892_ (
    .A(_00463_),
    .B(_00464_),
    .X(_00465_)
  );
  sg13g2_nor2_1 _10893_ (
    .A(_02294_),
    .B(_00465_),
    .Y(_00466_)
  );
  sg13g2_buf_1 _10894_ (
    .A(_00030_),
    .X(_00467_)
  );
  sg13g2_nand3_1 _10895_ (
    .A(addr_i_5_),
    .B(_00467_),
    .C(_02536_),
    .Y(_00468_)
  );
  sg13g2_a21oi_1 _10896_ (
    .A1(_00466_),
    .A2(_00468_),
    .B1(addr_i_8_),
    .Y(_00469_)
  );
  sg13g2_nand2_1 _10897_ (
    .A(addr_i_3_),
    .B(_05424_),
    .Y(_00470_)
  );
  sg13g2_nand2b_1 _10898_ (
    .A_N(_01417_),
    .B(_00470_),
    .Y(_00471_)
  );
  sg13g2_nor2_1 _10899_ (
    .A(addr_i_3_),
    .B(_06485_),
    .Y(_00472_)
  );
  sg13g2_buf_1 _10900_ (
    .A(_00472_),
    .X(_00474_)
  );
  sg13g2_a21oi_1 _10901_ (
    .A1(addr_i_7_),
    .A2(_00471_),
    .B1(_00474_),
    .Y(_00475_)
  );
  sg13g2_buf_1 _10902_ (
    .A(_01603_),
    .X(_00476_)
  );
  sg13g2_buf_1 _10903_ (
    .A(_01976_),
    .X(_00477_)
  );
  sg13g2_o21ai_1 _10904_ (
    .A1(_01153_),
    .A2(_03676_),
    .B1(addr_i_3_),
    .Y(_00478_)
  );
  sg13g2_buf_1 _10905_ (
    .A(_09038_),
    .X(_00479_)
  );
  sg13g2_o21ai_1 _10906_ (
    .A1(_00454_),
    .A2(_00014_),
    .B1(_00479_),
    .Y(_00480_)
  );
  sg13g2_nand4_1 _10907_ (
    .A(_00476_),
    .B(_00477_),
    .C(_00478_),
    .D(_00480_),
    .Y(_00481_)
  );
  sg13g2_buf_1 _10908_ (
    .A(_04715_),
    .X(_00482_)
  );
  sg13g2_buf_1 _10909_ (
    .A(_09038_),
    .X(_00483_)
  );
  sg13g2_buf_1 _10910_ (
    .A(_00483_),
    .X(_00485_)
  );
  sg13g2_a21oi_1 _10911_ (
    .A1(_04296_),
    .A2(_00482_),
    .B1(_00485_),
    .Y(_00486_)
  );
  sg13g2_a22oi_1 _10912_ (
    .A1(addr_i_4_),
    .A2(_00481_),
    .B1(_00486_),
    .B2(_05600_),
    .Y(_00487_)
  );
  sg13g2_o21ai_1 _10913_ (
    .A1(addr_i_4_),
    .A2(_00475_),
    .B1(_00487_),
    .Y(_00488_)
  );
  sg13g2_nand3_1 _10914_ (
    .A(_00467_),
    .B(_00428_),
    .C(_05557_),
    .Y(_00489_)
  );
  sg13g2_nand2_1 _10915_ (
    .A(addr_i_8_),
    .B(_00489_),
    .Y(_00490_)
  );
  sg13g2_buf_1 _10916_ (
    .A(_02141_),
    .X(_00491_)
  );
  sg13g2_buf_1 _10917_ (
    .A(_00435_),
    .X(_00492_)
  );
  sg13g2_a21oi_1 _10918_ (
    .A1(_00064_),
    .A2(_02591_),
    .B1(addr_i_3_),
    .Y(_00493_)
  );
  sg13g2_nor2_1 _10919_ (
    .A(_05845_),
    .B(_01625_),
    .Y(_00494_)
  );
  sg13g2_nor4_1 _10920_ (
    .A(_00491_),
    .B(_00492_),
    .C(_00493_),
    .D(_00494_),
    .Y(_00496_)
  );
  sg13g2_buf_1 _10921_ (
    .A(_00293_),
    .X(_00497_)
  );
  sg13g2_buf_1 _10922_ (
    .A(_08941_),
    .X(_00498_)
  );
  sg13g2_nand2_1 _10923_ (
    .A(_00692_),
    .B(_00498_),
    .Y(_00499_)
  );
  sg13g2_buf_1 _10924_ (
    .A(_05501_),
    .X(_00500_)
  );
  sg13g2_a22oi_1 _10925_ (
    .A1(_00497_),
    .A2(_00499_),
    .B1(_00500_),
    .B2(_00230_),
    .Y(_00501_)
  );
  sg13g2_nand2_1 _10926_ (
    .A(addr_i_3_),
    .B(_00173_),
    .Y(_00502_)
  );
  sg13g2_nor2_1 _10927_ (
    .A(addr_i_3_),
    .B(_04318_),
    .Y(_00503_)
  );
  sg13g2_nor2_1 _10928_ (
    .A(_00226_),
    .B(_00503_),
    .Y(_00504_)
  );
  sg13g2_buf_1 _10929_ (
    .A(_00025_),
    .X(_00505_)
  );
  sg13g2_buf_1 _10930_ (
    .A(_00505_),
    .X(_00507_)
  );
  sg13g2_a21oi_1 _10931_ (
    .A1(_00502_),
    .A2(_00504_),
    .B1(_00507_),
    .Y(_00508_)
  );
  sg13g2_nor4_1 _10932_ (
    .A(_00490_),
    .B(_00496_),
    .C(_00501_),
    .D(_00508_),
    .Y(_00509_)
  );
  sg13g2_a22oi_1 _10933_ (
    .A1(_00469_),
    .A2(_00488_),
    .B1(addr_i_9_),
    .B2(_00509_),
    .Y(_00510_)
  );
  sg13g2_buf_1 _10934_ (
    .A(_03731_),
    .X(_00511_)
  );
  sg13g2_a22oi_1 _10935_ (
    .A1(addr_i_9_),
    .A2(_00461_),
    .B1(_00510_),
    .B2(_00511_),
    .Y(_00512_)
  );
  sg13g2_nand2_1 _10936_ (
    .A(_02996_),
    .B(addr_i_11_),
    .Y(_00513_)
  );
  sg13g2_nor2_1 _10937_ (
    .A(_07226_),
    .B(_02097_),
    .Y(_00514_)
  );
  sg13g2_nor2_1 _10938_ (
    .A(addr_i_3_),
    .B(_00514_),
    .Y(_00515_)
  );
  sg13g2_buf_1 _10939_ (
    .A(_01757_),
    .X(_00516_)
  );
  sg13g2_nor2_1 _10940_ (
    .A(_00034_),
    .B(_00516_),
    .Y(_00518_)
  );
  sg13g2_o21ai_1 _10941_ (
    .A1(_00515_),
    .A2(_00518_),
    .B1(addr_i_2_),
    .Y(_00519_)
  );
  sg13g2_buf_1 _10942_ (
    .A(_04418_),
    .X(_00520_)
  );
  sg13g2_buf_1 _10943_ (
    .A(_01724_),
    .X(_00521_)
  );
  sg13g2_buf_1 _10944_ (
    .A(_00521_),
    .X(_00522_)
  );
  sg13g2_nor2_1 _10945_ (
    .A(_00520_),
    .B(_00522_),
    .Y(_00523_)
  );
  sg13g2_nor2_1 _10946_ (
    .A(addr_i_7_),
    .B(_00523_),
    .Y(_00524_)
  );
  sg13g2_a22oi_1 _10947_ (
    .A1(addr_i_2_),
    .A2(_08930_),
    .B1(_09459_),
    .B2(_08155_),
    .Y(_00525_)
  );
  sg13g2_o21ai_1 _10948_ (
    .A1(_00945_),
    .A2(_00525_),
    .B1(addr_i_3_),
    .Y(_00526_)
  );
  sg13g2_nand3_1 _10949_ (
    .A(_00519_),
    .B(_00524_),
    .C(_00526_),
    .Y(_00527_)
  );
  sg13g2_buf_1 _10950_ (
    .A(_09061_),
    .X(_00529_)
  );
  sg13g2_nand3_1 _10951_ (
    .A(_00529_),
    .B(_00224_),
    .C(_08620_),
    .Y(_00530_)
  );
  sg13g2_buf_1 _10952_ (
    .A(_00333_),
    .X(_00531_)
  );
  sg13g2_nor2_1 _10953_ (
    .A(_00531_),
    .B(_02755_),
    .Y(_00532_)
  );
  sg13g2_nor2_1 _10954_ (
    .A(_08299_),
    .B(_05999_),
    .Y(_00533_)
  );
  sg13g2_buf_1 _10955_ (
    .A(_02108_),
    .X(_00534_)
  );
  sg13g2_buf_1 _10956_ (
    .A(_05269_),
    .X(_00535_)
  );
  sg13g2_nor2_1 _10957_ (
    .A(_00535_),
    .B(_05036_),
    .Y(_00536_)
  );
  sg13g2_o21ai_1 _10958_ (
    .A1(_00534_),
    .A2(_00536_),
    .B1(addr_i_4_),
    .Y(_00537_)
  );
  sg13g2_o21ai_1 _10959_ (
    .A1(addr_i_3_),
    .A2(_00533_),
    .B1(_00537_),
    .Y(_00538_)
  );
  sg13g2_o21ai_1 _10960_ (
    .A1(_00532_),
    .A2(_00538_),
    .B1(addr_i_7_),
    .Y(_00540_)
  );
  sg13g2_nand4_1 _10961_ (
    .A(_03259_),
    .B(_00527_),
    .C(_00530_),
    .D(_00540_),
    .Y(_00541_)
  );
  sg13g2_buf_1 _10962_ (
    .A(_08852_),
    .X(_00542_)
  );
  sg13g2_buf_1 _10963_ (
    .A(_00521_),
    .X(_00543_)
  );
  sg13g2_nand2_1 _10964_ (
    .A(addr_i_5_),
    .B(_00543_),
    .Y(_00544_)
  );
  sg13g2_nand2_1 _10965_ (
    .A(_05346_),
    .B(_07492_),
    .Y(_00545_)
  );
  sg13g2_o21ai_1 _10966_ (
    .A1(_00542_),
    .A2(_00544_),
    .B1(_00545_),
    .Y(_00546_)
  );
  sg13g2_buf_1 _10967_ (
    .A(_04904_),
    .X(_00547_)
  );
  sg13g2_buf_1 _10968_ (
    .A(_00547_),
    .X(_00548_)
  );
  sg13g2_buf_1 _10969_ (
    .A(_08564_),
    .X(_00549_)
  );
  sg13g2_nand2_1 _10970_ (
    .A(_00549_),
    .B(_08254_),
    .Y(_00551_)
  );
  sg13g2_nor2_1 _10971_ (
    .A(_00536_),
    .B(_00551_),
    .Y(_00552_)
  );
  sg13g2_o21ai_1 _10972_ (
    .A1(_00548_),
    .A2(_00552_),
    .B1(addr_i_8_),
    .Y(_00553_)
  );
  sg13g2_buf_1 _10973_ (
    .A(_00342_),
    .X(_00554_)
  );
  sg13g2_a21oi_1 _10974_ (
    .A1(_04162_),
    .A2(_00358_),
    .B1(_00554_),
    .Y(_00555_)
  );
  sg13g2_nor2_1 _10975_ (
    .A(_09359_),
    .B(_00555_),
    .Y(_00556_)
  );
  sg13g2_buf_1 _10976_ (
    .A(_02108_),
    .X(_00557_)
  );
  sg13g2_nor3_1 _10977_ (
    .A(addr_i_4_),
    .B(_00014_),
    .C(_00557_),
    .Y(_00558_)
  );
  sg13g2_nor2_1 _10978_ (
    .A(_07933_),
    .B(_03490_),
    .Y(_00559_)
  );
  sg13g2_o21ai_1 _10979_ (
    .A1(_00558_),
    .A2(_00559_),
    .B1(addr_i_3_),
    .Y(_00560_)
  );
  sg13g2_a21oi_1 _10980_ (
    .A1(_00556_),
    .A2(_00560_),
    .B1(addr_i_7_),
    .Y(_00562_)
  );
  sg13g2_a22oi_1 _10981_ (
    .A1(_00169_),
    .A2(_00546_),
    .B1(_00553_),
    .B2(_00562_),
    .Y(_00563_)
  );
  sg13g2_nor2_1 _10982_ (
    .A(_00396_),
    .B(_00563_),
    .Y(_00564_)
  );
  sg13g2_buf_1 _10983_ (
    .A(_00059_),
    .X(_00565_)
  );
  sg13g2_buf_1 _10984_ (
    .A(_06077_),
    .X(_00566_)
  );
  sg13g2_nand2_1 _10985_ (
    .A(addr_i_4_),
    .B(_04860_),
    .Y(_00567_)
  );
  sg13g2_nand2_1 _10986_ (
    .A(_00566_),
    .B(_00567_),
    .Y(_00568_)
  );
  sg13g2_nor2_1 _10987_ (
    .A(_03446_),
    .B(_08941_),
    .Y(_00569_)
  );
  sg13g2_a21oi_1 _10988_ (
    .A1(_00565_),
    .A2(_00568_),
    .B1(_00569_),
    .Y(_00570_)
  );
  sg13g2_buf_1 _10989_ (
    .A(_01241_),
    .X(_00571_)
  );
  sg13g2_buf_1 _10990_ (
    .A(_00571_),
    .X(_00573_)
  );
  sg13g2_nand2_1 _10991_ (
    .A(addr_i_6_),
    .B(_01636_),
    .Y(_00574_)
  );
  sg13g2_a221oi_1 _10992_ (
    .A1(addr_i_5_),
    .A2(_00573_),
    .B1(_00574_),
    .B2(addr_i_3_),
    .C1(addr_i_2_),
    .Y(_00575_)
  );
  sg13g2_a22oi_1 _10993_ (
    .A1(addr_i_2_),
    .A2(_00570_),
    .B1(_00575_),
    .B2(_00290_),
    .Y(_00576_)
  );
  sg13g2_xor2_1 _10994_ (
    .A(addr_i_4_),
    .B(addr_i_6_),
    .X(_00577_)
  );
  sg13g2_buf_1 _10995_ (
    .A(_00577_),
    .X(_00578_)
  );
  sg13g2_nor2_1 _10996_ (
    .A(addr_i_3_),
    .B(_00578_),
    .Y(_00579_)
  );
  sg13g2_o21ai_1 _10997_ (
    .A1(_00334_),
    .A2(_00579_),
    .B1(addr_i_2_),
    .Y(_00580_)
  );
  sg13g2_buf_1 _10998_ (
    .A(_00462_),
    .X(_00581_)
  );
  sg13g2_buf_1 _10999_ (
    .A(_00581_),
    .X(_00582_)
  );
  sg13g2_nand2_1 _11000_ (
    .A(addr_i_4_),
    .B(_01976_),
    .Y(_00584_)
  );
  sg13g2_nand2_1 _11001_ (
    .A(_00582_),
    .B(_00584_),
    .Y(_00585_)
  );
  sg13g2_buf_1 _11002_ (
    .A(_00681_),
    .X(_00586_)
  );
  sg13g2_nor2_1 _11003_ (
    .A(_00586_),
    .B(_01570_),
    .Y(_00587_)
  );
  sg13g2_buf_1 _11004_ (
    .A(_01011_),
    .X(_00588_)
  );
  sg13g2_a22oi_1 _11005_ (
    .A1(addr_i_3_),
    .A2(_00585_),
    .B1(_00587_),
    .B2(_00588_),
    .Y(_00589_)
  );
  sg13g2_o21ai_1 _11006_ (
    .A1(addr_i_6_),
    .A2(addr_i_5_),
    .B1(addr_i_2_),
    .Y(_00590_)
  );
  sg13g2_buf_1 _11007_ (
    .A(_00590_),
    .X(_00591_)
  );
  sg13g2_or2_1 _11008_ (
    .A(_05856_),
    .B(_00591_),
    .X(_00592_)
  );
  sg13g2_buf_1 _11009_ (
    .A(_05269_),
    .X(_00593_)
  );
  sg13g2_nand2_1 _11010_ (
    .A(_00593_),
    .B(_05966_),
    .Y(_00595_)
  );
  sg13g2_nand3_1 _11011_ (
    .A(addr_i_4_),
    .B(_00592_),
    .C(_00595_),
    .Y(_00596_)
  );
  sg13g2_buf_1 _11012_ (
    .A(_06541_),
    .X(_00597_)
  );
  sg13g2_nor3_1 _11013_ (
    .A(addr_i_3_),
    .B(_08896_),
    .C(_03172_),
    .Y(_00598_)
  );
  sg13g2_or3_1 _11014_ (
    .A(addr_i_4_),
    .B(_00597_),
    .C(_00598_),
    .X(_00599_)
  );
  sg13g2_buf_1 _11015_ (
    .A(_07591_),
    .X(_00600_)
  );
  sg13g2_a21oi_1 _11016_ (
    .A1(_00596_),
    .A2(_00599_),
    .B1(_00600_),
    .Y(_00601_)
  );
  sg13g2_a21oi_1 _11017_ (
    .A1(_00580_),
    .A2(_00589_),
    .B1(_00601_),
    .Y(_00602_)
  );
  sg13g2_nand2_1 _11018_ (
    .A(addr_i_3_),
    .B(_08763_),
    .Y(_00603_)
  );
  sg13g2_nand2_1 _11019_ (
    .A(_00358_),
    .B(_00603_),
    .Y(_00604_)
  );
  sg13g2_a22oi_1 _11020_ (
    .A1(addr_i_5_),
    .A2(_00604_),
    .B1(_06574_),
    .B2(_00659_),
    .Y(_00606_)
  );
  sg13g2_buf_1 _11021_ (
    .A(_02503_),
    .X(_00607_)
  );
  sg13g2_nor2_1 _11022_ (
    .A(addr_i_3_),
    .B(_00327_),
    .Y(_00608_)
  );
  sg13g2_nor3_1 _11023_ (
    .A(addr_i_4_),
    .B(_00607_),
    .C(_00608_),
    .Y(_00609_)
  );
  sg13g2_buf_1 _11024_ (
    .A(_04650_),
    .X(_00610_)
  );
  sg13g2_o21ai_1 _11025_ (
    .A1(_00606_),
    .A2(_00609_),
    .B1(_00610_),
    .Y(_00611_)
  );
  sg13g2_nand3b_1 _11026_ (
    .A_N(_00576_),
    .B(_00602_),
    .C(_00611_),
    .Y(_00612_)
  );
  sg13g2_a221oi_1 _11027_ (
    .A1(_00541_),
    .A2(_00564_),
    .B1(_00612_),
    .B2(_00397_),
    .C1(addr_i_10_),
    .Y(_00613_)
  );
  sg13g2_nor3_1 _11028_ (
    .A(_00512_),
    .B(_00513_),
    .C(_00613_),
    .Y(_00614_)
  );
  sg13g2_a21oi_1 _11029_ (
    .A1(_00313_),
    .A2(_00425_),
    .B1(_00614_),
    .Y(_00615_)
  );
  sg13g2_o21ai_1 _11030_ (
    .A1(_00167_),
    .A2(_00218_),
    .B1(_00615_),
    .Y(data_o_10_)
  );
  sg13g2_buf_1 _11031_ (
    .A(_06220_),
    .X(_00617_)
  );
  sg13g2_or3_1 _11032_ (
    .A(addr_i_2_),
    .B(addr_i_7_),
    .C(addr_i_6_),
    .X(_00618_)
  );
  sg13g2_nand2_1 _11033_ (
    .A(_07050_),
    .B(_00618_),
    .Y(_00619_)
  );
  sg13g2_nand2_1 _11034_ (
    .A(_07491_),
    .B(_05225_),
    .Y(_00620_)
  );
  sg13g2_o21ai_1 _11035_ (
    .A1(addr_i_6_),
    .A2(_06729_),
    .B1(addr_i_5_),
    .Y(_00621_)
  );
  sg13g2_a21oi_1 _11036_ (
    .A1(_00620_),
    .A2(_00621_),
    .B1(addr_i_4_),
    .Y(_00622_)
  );
  sg13g2_a22oi_1 _11037_ (
    .A1(_00617_),
    .A2(_00619_),
    .B1(_00622_),
    .B2(addr_i_3_),
    .Y(_00623_)
  );
  sg13g2_buf_1 _11038_ (
    .A(_08597_),
    .X(_00624_)
  );
  sg13g2_o21ai_1 _11039_ (
    .A1(_00624_),
    .A2(_00165_),
    .B1(_07658_),
    .Y(_00625_)
  );
  sg13g2_a21oi_1 _11040_ (
    .A1(_00404_),
    .A2(_00625_),
    .B1(addr_i_4_),
    .Y(_00627_)
  );
  sg13g2_a22oi_1 _11041_ (
    .A1(_00261_),
    .A2(_04505_),
    .B1(_00627_),
    .B2(_00485_),
    .Y(_00628_)
  );
  sg13g2_buf_1 _11042_ (
    .A(_06684_),
    .X(_00629_)
  );
  sg13g2_o21ai_1 _11043_ (
    .A1(_00623_),
    .A2(_00628_),
    .B1(_00629_),
    .Y(_00630_)
  );
  sg13g2_and3_1 _11044_ (
    .A(addr_i_2_),
    .B(addr_i_7_),
    .C(addr_i_5_),
    .X(_00631_)
  );
  sg13g2_buf_1 _11045_ (
    .A(_00631_),
    .X(_00632_)
  );
  sg13g2_nand2_1 _11046_ (
    .A(_00605_),
    .B(_00632_),
    .Y(_00633_)
  );
  sg13g2_o21ai_1 _11047_ (
    .A1(_05346_),
    .A2(_00583_),
    .B1(_09485_),
    .Y(_00634_)
  );
  sg13g2_nor2b_1 _11048_ (
    .A(addr_i_3_),
    .B_N(addr_i_7_),
    .Y(_00635_)
  );
  sg13g2_nand3_1 _11049_ (
    .A(_00260_),
    .B(_01581_),
    .C(_00635_),
    .Y(_00636_)
  );
  sg13g2_nand3_1 _11050_ (
    .A(addr_i_2_),
    .B(_09050_),
    .C(_01943_),
    .Y(_00638_)
  );
  sg13g2_nand4_1 _11051_ (
    .A(_00633_),
    .B(_00634_),
    .C(_00636_),
    .D(_00638_),
    .Y(_00639_)
  );
  sg13g2_nand2_1 _11052_ (
    .A(addr_i_4_),
    .B(_00639_),
    .Y(_00640_)
  );
  sg13g2_nor2_1 _11053_ (
    .A(_02196_),
    .B(_00547_),
    .Y(_00641_)
  );
  sg13g2_a21oi_1 _11054_ (
    .A1(_07326_),
    .A2(_03953_),
    .B1(_00333_),
    .Y(_00642_)
  );
  sg13g2_o21ai_1 _11055_ (
    .A1(_00641_),
    .A2(_00642_),
    .B1(_01131_),
    .Y(_00643_)
  );
  sg13g2_buf_1 _11056_ (
    .A(_05424_),
    .X(_00644_)
  );
  sg13g2_buf_1 _11057_ (
    .A(_00635_),
    .X(_00645_)
  );
  sg13g2_nand2_1 _11058_ (
    .A(_00644_),
    .B(_00645_),
    .Y(_00646_)
  );
  sg13g2_nand4_1 _11059_ (
    .A(addr_i_8_),
    .B(_00640_),
    .C(_00643_),
    .D(_00646_),
    .Y(_00647_)
  );
  sg13g2_nor2_1 _11060_ (
    .A(addr_i_3_),
    .B(_06298_),
    .Y(_00649_)
  );
  sg13g2_buf_1 _11061_ (
    .A(_04628_),
    .X(_00650_)
  );
  sg13g2_buf_1 _11062_ (
    .A(_00650_),
    .X(_00651_)
  );
  sg13g2_a221oi_1 _11063_ (
    .A1(addr_i_3_),
    .A2(_09484_),
    .B1(_00649_),
    .B2(_00651_),
    .C1(_07945_),
    .Y(_00652_)
  );
  sg13g2_a22oi_1 _11064_ (
    .A1(_00630_),
    .A2(_00647_),
    .B1(_00652_),
    .B2(addr_i_10_),
    .Y(_00653_)
  );
  sg13g2_nor2_1 _11065_ (
    .A(_09509_),
    .B(_00534_),
    .Y(_00654_)
  );
  sg13g2_nand2_1 _11066_ (
    .A(_00099_),
    .B(_02152_),
    .Y(_00655_)
  );
  sg13g2_nand2_1 _11067_ (
    .A(_09485_),
    .B(_02503_),
    .Y(_00656_)
  );
  sg13g2_nand2_1 _11068_ (
    .A(_00655_),
    .B(_00656_),
    .Y(_00657_)
  );
  sg13g2_nand2_1 _11069_ (
    .A(_00550_),
    .B(_00099_),
    .Y(_00658_)
  );
  sg13g2_nand2_1 _11070_ (
    .A(_01680_),
    .B(_06209_),
    .Y(_00660_)
  );
  sg13g2_a21oi_1 _11071_ (
    .A1(_00658_),
    .A2(_00660_),
    .B1(addr_i_3_),
    .Y(_00661_)
  );
  sg13g2_a22oi_1 _11072_ (
    .A1(addr_i_3_),
    .A2(_00654_),
    .B1(_00657_),
    .B2(_00661_),
    .Y(_00662_)
  );
  sg13g2_xnor2_1 _11073_ (
    .A(addr_i_6_),
    .B(addr_i_5_),
    .Y(_00663_)
  );
  sg13g2_buf_1 _11074_ (
    .A(_00663_),
    .X(_00664_)
  );
  sg13g2_buf_1 _11075_ (
    .A(_00664_),
    .X(_00665_)
  );
  sg13g2_buf_1 _11076_ (
    .A(_00665_),
    .X(_00666_)
  );
  sg13g2_nor2_1 _11077_ (
    .A(addr_i_3_),
    .B(_00406_),
    .Y(_00667_)
  );
  sg13g2_nand2_1 _11078_ (
    .A(_04151_),
    .B(_06563_),
    .Y(_00668_)
  );
  sg13g2_nand3b_1 _11079_ (
    .A_N(addr_i_4_),
    .B(addr_i_2_),
    .C(addr_i_6_),
    .Y(_00669_)
  );
  sg13g2_buf_1 _11080_ (
    .A(_00669_),
    .X(_00671_)
  );
  sg13g2_a21o_1 _11081_ (
    .A1(_08520_),
    .A2(_00671_),
    .B1(_02207_),
    .X(_00672_)
  );
  sg13g2_a21oi_1 _11082_ (
    .A1(_00668_),
    .A2(_00672_),
    .B1(addr_i_7_),
    .Y(_00673_)
  );
  sg13g2_a21oi_1 _11083_ (
    .A1(_00666_),
    .A2(_00667_),
    .B1(_00673_),
    .Y(_00674_)
  );
  sg13g2_o21ai_1 _11084_ (
    .A1(addr_i_2_),
    .A2(_00662_),
    .B1(_00674_),
    .Y(_00675_)
  );
  sg13g2_buf_1 _11085_ (
    .A(_00000_),
    .X(_00676_)
  );
  sg13g2_nand2_1 _11086_ (
    .A(_00110_),
    .B(_00676_),
    .Y(_00677_)
  );
  sg13g2_nand2b_1 _11087_ (
    .A_N(addr_i_7_),
    .B(addr_i_5_),
    .Y(_00678_)
  );
  sg13g2_buf_1 _11088_ (
    .A(_00678_),
    .X(_00679_)
  );
  sg13g2_nand3b_1 _11089_ (
    .A_N(addr_i_5_),
    .B(addr_i_7_),
    .C(addr_i_2_),
    .Y(_00680_)
  );
  sg13g2_o21ai_1 _11090_ (
    .A1(_00679_),
    .A2(_00406_),
    .B1(_00680_),
    .Y(_00682_)
  );
  sg13g2_nor3_1 _11091_ (
    .A(addr_i_4_),
    .B(_08885_),
    .C(_00154_),
    .Y(_00683_)
  );
  sg13g2_o21ai_1 _11092_ (
    .A1(_00682_),
    .A2(_00683_),
    .B1(_06607_),
    .Y(_00684_)
  );
  sg13g2_and2_1 _11093_ (
    .A(_00677_),
    .B(_00684_),
    .X(_00685_)
  );
  sg13g2_o21ai_1 _11094_ (
    .A1(addr_i_6_),
    .A2(_04804_),
    .B1(_07160_),
    .Y(_00686_)
  );
  sg13g2_buf_1 _11095_ (
    .A(_07469_),
    .X(_00687_)
  );
  sg13g2_buf_1 _11096_ (
    .A(_01636_),
    .X(_00688_)
  );
  sg13g2_a21oi_1 _11097_ (
    .A1(_04396_),
    .A2(_00687_),
    .B1(_00688_),
    .Y(_00689_)
  );
  sg13g2_a22oi_1 _11098_ (
    .A1(_00268_),
    .A2(_00686_),
    .B1(_00689_),
    .B2(addr_i_3_),
    .Y(_00690_)
  );
  sg13g2_a22oi_1 _11099_ (
    .A1(addr_i_3_),
    .A2(_00685_),
    .B1(_00690_),
    .B2(addr_i_8_),
    .Y(_00691_)
  );
  sg13g2_a22oi_1 _11100_ (
    .A1(addr_i_8_),
    .A2(_00675_),
    .B1(_00691_),
    .B2(_03731_),
    .Y(_00693_)
  );
  sg13g2_o21ai_1 _11101_ (
    .A1(_00653_),
    .A2(_00693_),
    .B1(addr_i_9_),
    .Y(_00694_)
  );
  sg13g2_buf_1 _11102_ (
    .A(_05910_),
    .X(_00695_)
  );
  sg13g2_nand3_1 _11103_ (
    .A(addr_i_5_),
    .B(_00695_),
    .C(_00594_),
    .Y(_00696_)
  );
  sg13g2_buf_1 _11104_ (
    .A(_00586_),
    .X(_00697_)
  );
  sg13g2_nand3_1 _11105_ (
    .A(addr_i_6_),
    .B(_00697_),
    .C(_03853_),
    .Y(_00698_)
  );
  sg13g2_nand2_1 _11106_ (
    .A(_00696_),
    .B(_00698_),
    .Y(_00699_)
  );
  sg13g2_buf_1 _11107_ (
    .A(_05324_),
    .X(_00700_)
  );
  sg13g2_buf_1 _11108_ (
    .A(_00700_),
    .X(_00701_)
  );
  sg13g2_nand2_1 _11109_ (
    .A(_06275_),
    .B(_00714_),
    .Y(_00702_)
  );
  sg13g2_buf_1 _11110_ (
    .A(_01087_),
    .X(_00704_)
  );
  sg13g2_o21ai_1 _11111_ (
    .A1(_00343_),
    .A2(_00702_),
    .B1(_00704_),
    .Y(_00705_)
  );
  sg13g2_and2_1 _11112_ (
    .A(_00701_),
    .B(_00705_),
    .X(_00706_)
  );
  sg13g2_o21ai_1 _11113_ (
    .A1(_00699_),
    .A2(_00706_),
    .B1(_00440_),
    .Y(_00707_)
  );
  sg13g2_buf_1 _11114_ (
    .A(_07934_),
    .X(_00708_)
  );
  sg13g2_nor2_1 _11115_ (
    .A(_06795_),
    .B(_06497_),
    .Y(_00709_)
  );
  sg13g2_o21ai_1 _11116_ (
    .A1(addr_i_4_),
    .A2(_00709_),
    .B1(_06585_),
    .Y(_00710_)
  );
  sg13g2_xnor2_1 _11117_ (
    .A(addr_i_3_),
    .B(addr_i_2_),
    .Y(_00711_)
  );
  sg13g2_buf_1 _11118_ (
    .A(_00711_),
    .X(_00712_)
  );
  sg13g2_and2_1 _11119_ (
    .A(addr_i_8_),
    .B(addr_i_7_),
    .X(_00713_)
  );
  sg13g2_nand2_1 _11120_ (
    .A(_06496_),
    .B(_00713_),
    .Y(_00715_)
  );
  sg13g2_buf_1 _11121_ (
    .A(_05678_),
    .X(_00716_)
  );
  sg13g2_nor2_1 _11122_ (
    .A(_00715_),
    .B(_00716_),
    .Y(_00717_)
  );
  sg13g2_nand2b_1 _11123_ (
    .A_N(addr_i_3_),
    .B(addr_i_5_),
    .Y(_00718_)
  );
  sg13g2_buf_1 _11124_ (
    .A(_00718_),
    .X(_00719_)
  );
  sg13g2_nand3_1 _11125_ (
    .A(addr_i_6_),
    .B(_06851_),
    .C(_02503_),
    .Y(_00720_)
  );
  sg13g2_nor2_1 _11126_ (
    .A(_00044_),
    .B(_07469_),
    .Y(_00721_)
  );
  sg13g2_a22oi_1 _11127_ (
    .A1(_00719_),
    .A2(_00720_),
    .B1(_00721_),
    .B2(_01011_),
    .Y(_00722_)
  );
  sg13g2_a22oi_1 _11128_ (
    .A1(_00712_),
    .A2(_00717_),
    .B1(_00722_),
    .B2(_03073_),
    .Y(_00723_)
  );
  sg13g2_inv_1 _11129_ (
    .A(_00723_),
    .Y(_00724_)
  );
  sg13g2_buf_1 _11130_ (
    .A(_00463_),
    .X(_00726_)
  );
  sg13g2_nor2_1 _11131_ (
    .A(_07237_),
    .B(_03194_),
    .Y(_00727_)
  );
  sg13g2_o21ai_1 _11132_ (
    .A1(_00726_),
    .A2(_00727_),
    .B1(_01230_),
    .Y(_00728_)
  );
  sg13g2_nor2_1 _11133_ (
    .A(_04539_),
    .B(_07359_),
    .Y(_00729_)
  );
  sg13g2_o21ai_1 _11134_ (
    .A1(addr_i_5_),
    .A2(_00729_),
    .B1(_00276_),
    .Y(_00730_)
  );
  sg13g2_buf_1 _11135_ (
    .A(_02185_),
    .X(_00731_)
  );
  sg13g2_nor2_1 _11136_ (
    .A(_00731_),
    .B(_06398_),
    .Y(_00732_)
  );
  sg13g2_a22oi_1 _11137_ (
    .A1(_00388_),
    .A2(_00728_),
    .B1(_00730_),
    .B2(_00732_),
    .Y(_00733_)
  );
  sg13g2_a22oi_1 _11138_ (
    .A1(_00708_),
    .A2(_00710_),
    .B1(_00724_),
    .B2(_00733_),
    .Y(_00734_)
  );
  sg13g2_o21ai_1 _11139_ (
    .A1(_08100_),
    .A2(_01570_),
    .B1(_01658_),
    .Y(_00735_)
  );
  sg13g2_nand3_1 _11140_ (
    .A(addr_i_5_),
    .B(_09393_),
    .C(_08719_),
    .Y(_00737_)
  );
  sg13g2_nor2_1 _11141_ (
    .A(addr_i_3_),
    .B(addr_i_5_),
    .Y(_00738_)
  );
  sg13g2_nand2_1 _11142_ (
    .A(_04749_),
    .B(_00738_),
    .Y(_00739_)
  );
  sg13g2_a21oi_1 _11143_ (
    .A1(_00737_),
    .A2(_00739_),
    .B1(_02064_),
    .Y(_00740_)
  );
  sg13g2_a21oi_1 _11144_ (
    .A1(addr_i_3_),
    .A2(_00735_),
    .B1(_00740_),
    .Y(_00741_)
  );
  sg13g2_and3_1 _11145_ (
    .A(addr_i_2_),
    .B(addr_i_6_),
    .C(addr_i_5_),
    .X(_00742_)
  );
  sg13g2_buf_1 _11146_ (
    .A(_00742_),
    .X(_00743_)
  );
  sg13g2_buf_1 _11147_ (
    .A(_00637_),
    .X(_00744_)
  );
  sg13g2_mux2_1 _11148_ (
    .A0(addr_i_2_),
    .A1(addr_i_5_),
    .S(addr_i_6_),
    .X(_00745_)
  );
  sg13g2_nor3_1 _11149_ (
    .A(addr_i_3_),
    .B(addr_i_6_),
    .C(addr_i_5_),
    .Y(_00746_)
  );
  sg13g2_a21oi_1 _11150_ (
    .A1(addr_i_3_),
    .A2(_00745_),
    .B1(_00746_),
    .Y(_00748_)
  );
  sg13g2_nand2_1 _11151_ (
    .A(_05700_),
    .B(_00890_),
    .Y(_00749_)
  );
  sg13g2_o21ai_1 _11152_ (
    .A1(_00744_),
    .A2(_00748_),
    .B1(_00749_),
    .Y(_00750_)
  );
  sg13g2_a221oi_1 _11153_ (
    .A1(_00743_),
    .A2(_00522_),
    .B1(_00750_),
    .B2(addr_i_7_),
    .C1(addr_i_8_),
    .Y(_00751_)
  );
  sg13g2_o21ai_1 _11154_ (
    .A1(addr_i_4_),
    .A2(_00741_),
    .B1(_00751_),
    .Y(_00752_)
  );
  sg13g2_a21oi_1 _11155_ (
    .A1(_04063_),
    .A2(_00477_),
    .B1(_00046_),
    .Y(_00753_)
  );
  sg13g2_nand2_1 _11156_ (
    .A(addr_i_5_),
    .B(_00327_),
    .Y(_00754_)
  );
  sg13g2_nor2_1 _11157_ (
    .A(_02602_),
    .B(_06574_),
    .Y(_00755_)
  );
  sg13g2_a21oi_1 _11158_ (
    .A1(addr_i_4_),
    .A2(_00754_),
    .B1(_00755_),
    .Y(_00756_)
  );
  sg13g2_o21ai_1 _11159_ (
    .A1(_00753_),
    .A2(_00756_),
    .B1(addr_i_7_),
    .Y(_00757_)
  );
  sg13g2_a21oi_1 _11160_ (
    .A1(addr_i_7_),
    .A2(addr_i_5_),
    .B1(addr_i_2_),
    .Y(_00759_)
  );
  sg13g2_nor2_1 _11161_ (
    .A(_00454_),
    .B(_00759_),
    .Y(_00760_)
  );
  sg13g2_nor2_1 _11162_ (
    .A(_05745_),
    .B(_00760_),
    .Y(_00761_)
  );
  sg13g2_nand2_1 _11163_ (
    .A(addr_i_3_),
    .B(_08885_),
    .Y(_00762_)
  );
  sg13g2_nand3b_1 _11164_ (
    .A_N(addr_i_7_),
    .B(addr_i_5_),
    .C(addr_i_2_),
    .Y(_00763_)
  );
  sg13g2_buf_1 _11165_ (
    .A(_00763_),
    .X(_00764_)
  );
  sg13g2_a21oi_1 _11166_ (
    .A1(_00762_),
    .A2(_00764_),
    .B1(addr_i_4_),
    .Y(_00765_)
  );
  sg13g2_o21ai_1 _11167_ (
    .A1(_00761_),
    .A2(_00765_),
    .B1(addr_i_6_),
    .Y(_00766_)
  );
  sg13g2_nand3_1 _11168_ (
    .A(addr_i_8_),
    .B(_00757_),
    .C(_00766_),
    .Y(_00767_)
  );
  sg13g2_xor2_1 _11169_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .X(_00768_)
  );
  sg13g2_buf_1 _11170_ (
    .A(_00768_),
    .X(_00770_)
  );
  sg13g2_nand2_1 _11171_ (
    .A(addr_i_3_),
    .B(_00770_),
    .Y(_00771_)
  );
  sg13g2_a22oi_1 _11172_ (
    .A1(_00224_),
    .A2(_00771_),
    .B1(_00290_),
    .B2(_00403_),
    .Y(_00772_)
  );
  sg13g2_nor2_1 _11173_ (
    .A(addr_i_10_),
    .B(addr_i_9_),
    .Y(_00773_)
  );
  sg13g2_inv_1 _11174_ (
    .A(_00773_),
    .Y(_00774_)
  );
  sg13g2_a22oi_1 _11175_ (
    .A1(_00752_),
    .A2(_00767_),
    .B1(_00772_),
    .B2(_00774_),
    .Y(_00775_)
  );
  sg13g2_a22oi_1 _11176_ (
    .A1(_00707_),
    .A2(_00734_),
    .B1(_00775_),
    .B2(addr_i_11_),
    .Y(_00776_)
  );
  sg13g2_nand2_1 _11177_ (
    .A(_00694_),
    .B(_00776_),
    .Y(_00777_)
  );
  sg13g2_buf_1 _11178_ (
    .A(_03809_),
    .X(_00778_)
  );
  sg13g2_buf_1 _11179_ (
    .A(_00778_),
    .X(_00779_)
  );
  sg13g2_a22oi_1 _11180_ (
    .A1(addr_i_8_),
    .A2(_08774_),
    .B1(_00779_),
    .B2(_02700_),
    .Y(_00781_)
  );
  sg13g2_buf_1 _11181_ (
    .A(_00112_),
    .X(_00782_)
  );
  sg13g2_buf_1 _11182_ (
    .A(_00210_),
    .X(_00783_)
  );
  sg13g2_nand3b_1 _11183_ (
    .A_N(addr_i_4_),
    .B(addr_i_6_),
    .C(addr_i_5_),
    .Y(_00784_)
  );
  sg13g2_buf_1 _11184_ (
    .A(_00784_),
    .X(_00785_)
  );
  sg13g2_nand2_1 _11185_ (
    .A(_00198_),
    .B(_00785_),
    .Y(_00786_)
  );
  sg13g2_nor3_1 _11186_ (
    .A(addr_i_6_),
    .B(_06862_),
    .C(_02503_),
    .Y(_00787_)
  );
  sg13g2_a21oi_1 _11187_ (
    .A1(_00783_),
    .A2(_00786_),
    .B1(_00787_),
    .Y(_00788_)
  );
  sg13g2_nand2b_1 _11188_ (
    .A_N(addr_i_7_),
    .B(addr_i_3_),
    .Y(_00789_)
  );
  sg13g2_a21oi_1 _11189_ (
    .A1(_03676_),
    .A2(_00789_),
    .B1(_05966_),
    .Y(_00790_)
  );
  sg13g2_nor2_1 _11190_ (
    .A(addr_i_3_),
    .B(_00246_),
    .Y(_00792_)
  );
  sg13g2_nor4_1 _11191_ (
    .A(_00086_),
    .B(_08852_),
    .C(_00790_),
    .D(_00792_),
    .Y(_00793_)
  );
  sg13g2_nor2_1 _11192_ (
    .A(_09415_),
    .B(_00543_),
    .Y(_00794_)
  );
  sg13g2_a21oi_1 _11193_ (
    .A1(addr_i_4_),
    .A2(_00793_),
    .B1(_00794_),
    .Y(_00795_)
  );
  sg13g2_o21ai_1 _11194_ (
    .A1(addr_i_7_),
    .A2(_00788_),
    .B1(_00795_),
    .Y(_00796_)
  );
  sg13g2_nand2_1 _11195_ (
    .A(_06364_),
    .B(_05678_),
    .Y(_00797_)
  );
  sg13g2_nor2_1 _11196_ (
    .A(_03919_),
    .B(_00797_),
    .Y(_00798_)
  );
  sg13g2_buf_1 _11197_ (
    .A(_08785_),
    .X(_00799_)
  );
  sg13g2_o21ai_1 _11198_ (
    .A1(_07425_),
    .A2(_00798_),
    .B1(_00799_),
    .Y(_00800_)
  );
  sg13g2_nand2_1 _11199_ (
    .A(_02503_),
    .B(_00447_),
    .Y(_00801_)
  );
  sg13g2_a21o_1 _11200_ (
    .A1(_01768_),
    .A2(_00801_),
    .B1(addr_i_4_),
    .X(_00803_)
  );
  sg13g2_a21oi_1 _11201_ (
    .A1(_00800_),
    .A2(_00803_),
    .B1(_08674_),
    .Y(_00804_)
  );
  sg13g2_a22oi_1 _11202_ (
    .A1(_00782_),
    .A2(_00796_),
    .B1(_00804_),
    .B2(addr_i_9_),
    .Y(_00805_)
  );
  sg13g2_nor3_1 _11203_ (
    .A(addr_i_10_),
    .B(_00781_),
    .C(_00805_),
    .Y(_00806_)
  );
  sg13g2_nand2_1 _11204_ (
    .A(addr_i_10_),
    .B(_00422_),
    .Y(_00807_)
  );
  sg13g2_nor2_1 _11205_ (
    .A(addr_i_7_),
    .B(_00447_),
    .Y(_00808_)
  );
  sg13g2_a21oi_1 _11206_ (
    .A1(_04439_),
    .A2(_07911_),
    .B1(_00808_),
    .Y(_00809_)
  );
  sg13g2_nor2_1 _11207_ (
    .A(_00807_),
    .B(_00809_),
    .Y(_00810_)
  );
  sg13g2_o21ai_1 _11208_ (
    .A1(_00806_),
    .A2(_00810_),
    .B1(addr_i_11_),
    .Y(_00811_)
  );
  sg13g2_buf_1 _11209_ (
    .A(_02996_),
    .X(_00812_)
  );
  sg13g2_a21oi_1 _11210_ (
    .A1(_00777_),
    .A2(_00811_),
    .B1(_00812_),
    .Y(_00814_)
  );
  sg13g2_nand2_1 _11211_ (
    .A(_03776_),
    .B(_02525_),
    .Y(_00815_)
  );
  sg13g2_o21ai_1 _11212_ (
    .A1(_07746_),
    .A2(_09083_),
    .B1(addr_i_3_),
    .Y(_00816_)
  );
  sg13g2_o21ai_1 _11213_ (
    .A1(addr_i_3_),
    .A2(_00815_),
    .B1(_00816_),
    .Y(_00817_)
  );
  sg13g2_buf_1 _11214_ (
    .A(_01472_),
    .X(_00818_)
  );
  sg13g2_buf_1 _11215_ (
    .A(_00718_),
    .X(_00819_)
  );
  sg13g2_buf_1 _11216_ (
    .A(_00819_),
    .X(_00820_)
  );
  sg13g2_nand2_1 _11217_ (
    .A(_00818_),
    .B(_00820_),
    .Y(_00821_)
  );
  sg13g2_buf_1 _11218_ (
    .A(_00463_),
    .X(_00822_)
  );
  sg13g2_o21ai_1 _11219_ (
    .A1(_00415_),
    .A2(_00177_),
    .B1(_00822_),
    .Y(_00823_)
  );
  sg13g2_buf_1 _11220_ (
    .A(_00052_),
    .X(_00825_)
  );
  sg13g2_a21oi_1 _11221_ (
    .A1(_00821_),
    .A2(_00823_),
    .B1(_00825_),
    .Y(_00826_)
  );
  sg13g2_buf_1 _11222_ (
    .A(_06298_),
    .X(_00827_)
  );
  sg13g2_nor2_1 _11223_ (
    .A(_03369_),
    .B(_02645_),
    .Y(_00828_)
  );
  sg13g2_nor2_1 _11224_ (
    .A(_07326_),
    .B(_00828_),
    .Y(_00829_)
  );
  sg13g2_o21ai_1 _11225_ (
    .A1(_00827_),
    .A2(_00829_),
    .B1(_01878_),
    .Y(_00830_)
  );
  sg13g2_buf_1 _11226_ (
    .A(_04628_),
    .X(_00831_)
  );
  sg13g2_nand2_1 _11227_ (
    .A(_05269_),
    .B(_02525_),
    .Y(_00832_)
  );
  sg13g2_nand3_1 _11228_ (
    .A(_00831_),
    .B(_00314_),
    .C(_00832_),
    .Y(_00833_)
  );
  sg13g2_a21oi_1 _11229_ (
    .A1(_05247_),
    .A2(_00833_),
    .B1(_05888_),
    .Y(_00834_)
  );
  sg13g2_nand2_1 _11230_ (
    .A(_00830_),
    .B(_00834_),
    .Y(_00836_)
  );
  sg13g2_a22oi_1 _11231_ (
    .A1(_00529_),
    .A2(_00817_),
    .B1(_00826_),
    .B2(_00836_),
    .Y(_00837_)
  );
  sg13g2_buf_1 _11232_ (
    .A(_03106_),
    .X(_00838_)
  );
  sg13g2_nor2_1 _11233_ (
    .A(addr_i_3_),
    .B(_03303_),
    .Y(_00839_)
  );
  sg13g2_buf_1 _11234_ (
    .A(_04086_),
    .X(_00840_)
  );
  sg13g2_o21ai_1 _11235_ (
    .A1(_00838_),
    .A2(_00839_),
    .B1(_00840_),
    .Y(_00841_)
  );
  sg13g2_nor2_1 _11236_ (
    .A(addr_i_5_),
    .B(_00578_),
    .Y(_00842_)
  );
  sg13g2_nand2_1 _11237_ (
    .A(_00322_),
    .B(_00842_),
    .Y(_00843_)
  );
  sg13g2_buf_1 _11238_ (
    .A(_08863_),
    .X(_00844_)
  );
  sg13g2_nand2_1 _11239_ (
    .A(_00783_),
    .B(_00844_),
    .Y(_00845_)
  );
  sg13g2_nand3_1 _11240_ (
    .A(_00841_),
    .B(_00843_),
    .C(_00845_),
    .Y(_00847_)
  );
  sg13g2_nand2_1 _11241_ (
    .A(_06862_),
    .B(_00650_),
    .Y(_00848_)
  );
  sg13g2_nand2_1 _11242_ (
    .A(_05867_),
    .B(_00848_),
    .Y(_00849_)
  );
  sg13g2_nor2_1 _11243_ (
    .A(_01373_),
    .B(_02722_),
    .Y(_00850_)
  );
  sg13g2_nor2_1 _11244_ (
    .A(_06375_),
    .B(_00850_),
    .Y(_00851_)
  );
  sg13g2_nand2_1 _11245_ (
    .A(addr_i_3_),
    .B(_07956_),
    .Y(_00852_)
  );
  sg13g2_nand2_1 _11246_ (
    .A(_00408_),
    .B(_00852_),
    .Y(_00853_)
  );
  sg13g2_nor3_1 _11247_ (
    .A(_04108_),
    .B(addr_i_2_),
    .C(_01954_),
    .Y(_00854_)
  );
  sg13g2_a22oi_1 _11248_ (
    .A1(addr_i_5_),
    .A2(_00853_),
    .B1(_00854_),
    .B2(addr_i_6_),
    .Y(_00855_)
  );
  sg13g2_a22oi_1 _11249_ (
    .A1(_00849_),
    .A2(_00851_),
    .B1(addr_i_7_),
    .B2(_00855_),
    .Y(_00856_)
  );
  sg13g2_a22oi_1 _11250_ (
    .A1(addr_i_7_),
    .A2(_00847_),
    .B1(_00856_),
    .B2(addr_i_8_),
    .Y(_00858_)
  );
  sg13g2_o21ai_1 _11251_ (
    .A1(_00837_),
    .A2(_00858_),
    .B1(addr_i_9_),
    .Y(_00859_)
  );
  sg13g2_buf_1 _11252_ (
    .A(_07591_),
    .X(_00860_)
  );
  sg13g2_buf_1 _11253_ (
    .A(_00583_),
    .X(_00861_)
  );
  sg13g2_nand2_1 _11254_ (
    .A(_08796_),
    .B(_00147_),
    .Y(_00862_)
  );
  sg13g2_nand2_1 _11255_ (
    .A(_00033_),
    .B(_02097_),
    .Y(_00863_)
  );
  sg13g2_nand2_1 _11256_ (
    .A(_00539_),
    .B(_01461_),
    .Y(_00864_)
  );
  sg13g2_a21oi_1 _11257_ (
    .A1(_00863_),
    .A2(_00864_),
    .B1(addr_i_3_),
    .Y(_00865_)
  );
  sg13g2_nor2_1 _11258_ (
    .A(_01965_),
    .B(_00521_),
    .Y(_00866_)
  );
  sg13g2_a22oi_1 _11259_ (
    .A1(_00861_),
    .A2(_00862_),
    .B1(_00865_),
    .B2(_00866_),
    .Y(_00867_)
  );
  sg13g2_or3_1 _11260_ (
    .A(addr_i_3_),
    .B(addr_i_2_),
    .C(addr_i_5_),
    .X(_00869_)
  );
  sg13g2_buf_1 _11261_ (
    .A(_00869_),
    .X(_00870_)
  );
  sg13g2_nand2_1 _11262_ (
    .A(_07933_),
    .B(_00495_),
    .Y(_00871_)
  );
  sg13g2_nand2_1 _11263_ (
    .A(_05335_),
    .B(_07447_),
    .Y(_00872_)
  );
  sg13g2_nand2_1 _11264_ (
    .A(_05269_),
    .B(_01625_),
    .Y(_00873_)
  );
  sg13g2_nand3_1 _11265_ (
    .A(_00871_),
    .B(_00872_),
    .C(_00873_),
    .Y(_00874_)
  );
  sg13g2_a221oi_1 _11266_ (
    .A1(_03380_),
    .A2(_00590_),
    .B1(_00874_),
    .B2(addr_i_6_),
    .C1(_00399_),
    .Y(_00875_)
  );
  sg13g2_a21o_1 _11267_ (
    .A1(_00870_),
    .A2(_00875_),
    .B1(_01494_),
    .X(_00876_)
  );
  sg13g2_o21ai_1 _11268_ (
    .A1(_00860_),
    .A2(_00867_),
    .B1(_00876_),
    .Y(_00877_)
  );
  sg13g2_buf_1 _11269_ (
    .A(_01987_),
    .X(_00878_)
  );
  sg13g2_o21ai_1 _11270_ (
    .A1(_00571_),
    .A2(_02755_),
    .B1(_00878_),
    .Y(_00880_)
  );
  sg13g2_a21oi_1 _11271_ (
    .A1(addr_i_3_),
    .A2(_00880_),
    .B1(_00399_),
    .Y(_00881_)
  );
  sg13g2_nor2_1 _11272_ (
    .A(_08830_),
    .B(_00881_),
    .Y(_00882_)
  );
  sg13g2_nand2_1 _11273_ (
    .A(addr_i_3_),
    .B(_08863_),
    .Y(_00883_)
  );
  sg13g2_buf_1 _11274_ (
    .A(_00883_),
    .X(_00884_)
  );
  sg13g2_nor2_1 _11275_ (
    .A(addr_i_3_),
    .B(_04793_),
    .Y(_00885_)
  );
  sg13g2_nor2_1 _11276_ (
    .A(addr_i_2_),
    .B(_00885_),
    .Y(_00886_)
  );
  sg13g2_nor2_1 _11277_ (
    .A(_00067_),
    .B(_00149_),
    .Y(_00887_)
  );
  sg13g2_a22oi_1 _11278_ (
    .A1(_00884_),
    .A2(_00886_),
    .B1(_00887_),
    .B2(_00588_),
    .Y(_00888_)
  );
  sg13g2_or4_1 _11279_ (
    .A(addr_i_9_),
    .B(_00877_),
    .C(_00882_),
    .D(_00888_),
    .X(_00889_)
  );
  sg13g2_nand3_1 _11280_ (
    .A(_00511_),
    .B(_00859_),
    .C(_00889_),
    .Y(_00891_)
  );
  sg13g2_o21ai_1 _11281_ (
    .A1(addr_i_6_),
    .A2(_00712_),
    .B1(_00200_),
    .Y(_00892_)
  );
  sg13g2_a21oi_1 _11282_ (
    .A1(_00737_),
    .A2(_00892_),
    .B1(addr_i_4_),
    .Y(_00893_)
  );
  sg13g2_nand2_1 _11283_ (
    .A(addr_i_3_),
    .B(_04749_),
    .Y(_00894_)
  );
  sg13g2_nand3_1 _11284_ (
    .A(addr_i_4_),
    .B(_00894_),
    .C(_00737_),
    .Y(_00895_)
  );
  sg13g2_nand2b_1 _11285_ (
    .A_N(_00893_),
    .B(_00895_),
    .Y(_00896_)
  );
  sg13g2_nor2_1 _11286_ (
    .A(addr_i_5_),
    .B(_04561_),
    .Y(_00897_)
  );
  sg13g2_buf_1 _11287_ (
    .A(_00897_),
    .X(_00898_)
  );
  sg13g2_buf_1 _11288_ (
    .A(_00505_),
    .X(_00899_)
  );
  sg13g2_nor3_1 _11289_ (
    .A(_00899_),
    .B(_02755_),
    .C(_00127_),
    .Y(_00900_)
  );
  sg13g2_a22oi_1 _11290_ (
    .A1(_00898_),
    .A2(_00853_),
    .B1(_00900_),
    .B2(addr_i_8_),
    .Y(_00902_)
  );
  sg13g2_o21ai_1 _11291_ (
    .A1(addr_i_7_),
    .A2(_00896_),
    .B1(_00902_),
    .Y(_00903_)
  );
  sg13g2_nand2_1 _11292_ (
    .A(_01581_),
    .B(_03314_),
    .Y(_00904_)
  );
  sg13g2_o21ai_1 _11293_ (
    .A1(addr_i_3_),
    .A2(_00904_),
    .B1(_02887_),
    .Y(_00905_)
  );
  sg13g2_nand2_1 _11294_ (
    .A(_00024_),
    .B(_03139_),
    .Y(_00906_)
  );
  sg13g2_nand2_1 _11295_ (
    .A(_04528_),
    .B(_06530_),
    .Y(_00907_)
  );
  sg13g2_a21oi_1 _11296_ (
    .A1(_00906_),
    .A2(_00907_),
    .B1(_02404_),
    .Y(_00908_)
  );
  sg13g2_a21o_1 _11297_ (
    .A1(addr_i_2_),
    .A2(_00905_),
    .B1(_00908_),
    .X(_00909_)
  );
  sg13g2_buf_1 _11298_ (
    .A(_00483_),
    .X(_00910_)
  );
  sg13g2_a21oi_1 _11299_ (
    .A1(_07491_),
    .A2(_02097_),
    .B1(_01142_),
    .Y(_00911_)
  );
  sg13g2_nand2_1 _11300_ (
    .A(_00910_),
    .B(_00911_),
    .Y(_00913_)
  );
  sg13g2_buf_1 _11301_ (
    .A(_01373_),
    .X(_00914_)
  );
  sg13g2_buf_1 _11302_ (
    .A(_00923_),
    .X(_00915_)
  );
  sg13g2_nand3_1 _11303_ (
    .A(addr_i_4_),
    .B(_00914_),
    .C(_00915_),
    .Y(_00916_)
  );
  sg13g2_nor2_1 _11304_ (
    .A(_00242_),
    .B(_01153_),
    .Y(_00917_)
  );
  sg13g2_nand2_1 _11305_ (
    .A(_00648_),
    .B(_00917_),
    .Y(_00918_)
  );
  sg13g2_nand3_1 _11306_ (
    .A(addr_i_3_),
    .B(_00916_),
    .C(_00918_),
    .Y(_00919_)
  );
  sg13g2_nor3_1 _11307_ (
    .A(addr_i_4_),
    .B(addr_i_6_),
    .C(_02503_),
    .Y(_00920_)
  );
  sg13g2_a22oi_1 _11308_ (
    .A1(_00913_),
    .A2(_00919_),
    .B1(_06905_),
    .B2(_00920_),
    .Y(_00921_)
  );
  sg13g2_a22oi_1 _11309_ (
    .A1(_06630_),
    .A2(_00909_),
    .B1(_00921_),
    .B2(_07293_),
    .Y(_00922_)
  );
  sg13g2_nor2_1 _11310_ (
    .A(_06652_),
    .B(_00922_),
    .Y(_00924_)
  );
  sg13g2_buf_1 _11311_ (
    .A(_00108_),
    .X(_00925_)
  );
  sg13g2_nand3b_1 _11312_ (
    .A_N(addr_i_7_),
    .B(addr_i_2_),
    .C(addr_i_4_),
    .Y(_00926_)
  );
  sg13g2_buf_1 _11313_ (
    .A(_06972_),
    .X(_00927_)
  );
  sg13g2_nand3_1 _11314_ (
    .A(_00927_),
    .B(_08930_),
    .C(_07967_),
    .Y(_00928_)
  );
  sg13g2_nand2_1 _11315_ (
    .A(_00926_),
    .B(_00928_),
    .Y(_00929_)
  );
  sg13g2_buf_1 _11316_ (
    .A(_04494_),
    .X(_00930_)
  );
  sg13g2_a21oi_1 _11317_ (
    .A1(_00692_),
    .A2(_08464_),
    .B1(_00930_),
    .Y(_00931_)
  );
  sg13g2_o21ai_1 _11318_ (
    .A1(_00667_),
    .A2(_00931_),
    .B1(addr_i_5_),
    .Y(_00932_)
  );
  sg13g2_nor2_1 _11319_ (
    .A(_00593_),
    .B(_06972_),
    .Y(_00933_)
  );
  sg13g2_a22oi_1 _11320_ (
    .A1(_00156_),
    .A2(_00302_),
    .B1(_00933_),
    .B2(_00017_),
    .Y(_00935_)
  );
  sg13g2_a21oi_1 _11321_ (
    .A1(_00932_),
    .A2(_00935_),
    .B1(addr_i_6_),
    .Y(_00936_)
  );
  sg13g2_a22oi_1 _11322_ (
    .A1(addr_i_3_),
    .A2(_00929_),
    .B1(_00936_),
    .B2(_07293_),
    .Y(_00937_)
  );
  sg13g2_buf_1 _11323_ (
    .A(_06485_),
    .X(_00938_)
  );
  sg13g2_nand2_1 _11324_ (
    .A(addr_i_2_),
    .B(_00938_),
    .Y(_00939_)
  );
  sg13g2_nand2_1 _11325_ (
    .A(_05269_),
    .B(_02909_),
    .Y(_00940_)
  );
  sg13g2_nand2_1 _11326_ (
    .A(_00137_),
    .B(_00940_),
    .Y(_00941_)
  );
  sg13g2_a21oi_1 _11327_ (
    .A1(addr_i_3_),
    .A2(_00939_),
    .B1(_00941_),
    .Y(_00942_)
  );
  sg13g2_nand2_1 _11328_ (
    .A(addr_i_3_),
    .B(_05966_),
    .Y(_00943_)
  );
  sg13g2_o21ai_1 _11329_ (
    .A1(_00659_),
    .A2(_00942_),
    .B1(_00943_),
    .Y(_00944_)
  );
  sg13g2_nor2_1 _11330_ (
    .A(_07381_),
    .B(_02272_),
    .Y(_00946_)
  );
  sg13g2_nor2_1 _11331_ (
    .A(_05281_),
    .B(_00413_),
    .Y(_00947_)
  );
  sg13g2_o21ai_1 _11332_ (
    .A1(_00946_),
    .A2(_00947_),
    .B1(addr_i_5_),
    .Y(_00948_)
  );
  sg13g2_buf_1 _11333_ (
    .A(_03776_),
    .X(_00949_)
  );
  sg13g2_nand2_1 _11334_ (
    .A(_07049_),
    .B(_03798_),
    .Y(_00950_)
  );
  sg13g2_buf_1 _11335_ (
    .A(_00950_),
    .X(_00951_)
  );
  sg13g2_o21ai_1 _11336_ (
    .A1(_00448_),
    .A2(_00951_),
    .B1(_08232_),
    .Y(_00952_)
  );
  sg13g2_nand2_1 _11337_ (
    .A(_00949_),
    .B(_00952_),
    .Y(_00953_)
  );
  sg13g2_a21oi_1 _11338_ (
    .A1(_00948_),
    .A2(_00953_),
    .B1(addr_i_4_),
    .Y(_00954_)
  );
  sg13g2_a22oi_1 _11339_ (
    .A1(addr_i_7_),
    .A2(_00944_),
    .B1(_00954_),
    .B2(addr_i_8_),
    .Y(_00955_)
  );
  sg13g2_nor3_1 _11340_ (
    .A(_00925_),
    .B(_00937_),
    .C(_00955_),
    .Y(_00957_)
  );
  sg13g2_a22oi_1 _11341_ (
    .A1(_00903_),
    .A2(_00924_),
    .B1(_03040_),
    .B2(_00957_),
    .Y(_00958_)
  );
  sg13g2_buf_1 _11342_ (
    .A(_08089_),
    .X(_00959_)
  );
  sg13g2_buf_1 _11343_ (
    .A(_07447_),
    .X(_00960_)
  );
  sg13g2_nand2b_1 _11344_ (
    .A_N(addr_i_3_),
    .B(addr_i_7_),
    .Y(_00961_)
  );
  sg13g2_a21oi_1 _11345_ (
    .A1(_06132_),
    .A2(_00671_),
    .B1(_00961_),
    .Y(_00962_)
  );
  sg13g2_a221oi_1 _11346_ (
    .A1(addr_i_4_),
    .A2(_00959_),
    .B1(_00100_),
    .B2(_00960_),
    .C1(_00962_),
    .Y(_00963_)
  );
  sg13g2_or2_1 _11347_ (
    .A(addr_i_4_),
    .B(addr_i_7_),
    .X(_00964_)
  );
  sg13g2_buf_1 _11348_ (
    .A(_00964_),
    .X(_00965_)
  );
  sg13g2_nand2_1 _11349_ (
    .A(_00549_),
    .B(_00965_),
    .Y(_00966_)
  );
  sg13g2_nand2_1 _11350_ (
    .A(_00120_),
    .B(_00006_),
    .Y(_00968_)
  );
  sg13g2_nor2_1 _11351_ (
    .A(addr_i_4_),
    .B(_00968_),
    .Y(_00969_)
  );
  sg13g2_a22oi_1 _11352_ (
    .A1(_01450_),
    .A2(_00966_),
    .B1(_00969_),
    .B2(addr_i_5_),
    .Y(_00970_)
  );
  sg13g2_a21oi_1 _11353_ (
    .A1(addr_i_5_),
    .A2(_00963_),
    .B1(_00970_),
    .Y(_00971_)
  );
  sg13g2_buf_1 _11354_ (
    .A(_00008_),
    .X(_00972_)
  );
  sg13g2_nand3b_1 _11355_ (
    .A_N(addr_i_2_),
    .B(addr_i_7_),
    .C(addr_i_3_),
    .Y(_00973_)
  );
  sg13g2_nand2_1 _11356_ (
    .A(_00731_),
    .B(_00973_),
    .Y(_00974_)
  );
  sg13g2_nand3b_1 _11357_ (
    .A_N(addr_i_2_),
    .B(addr_i_7_),
    .C(addr_i_4_),
    .Y(_00975_)
  );
  sg13g2_a21oi_1 _11358_ (
    .A1(_00965_),
    .A2(_00975_),
    .B1(_00819_),
    .Y(_00976_)
  );
  sg13g2_nor2_1 _11359_ (
    .A(addr_i_5_),
    .B(_04804_),
    .Y(_00977_)
  );
  sg13g2_a22oi_1 _11360_ (
    .A1(_00972_),
    .A2(_00974_),
    .B1(_00976_),
    .B2(_00977_),
    .Y(_00979_)
  );
  sg13g2_nand2_1 _11361_ (
    .A(_07061_),
    .B(_00557_),
    .Y(_00980_)
  );
  sg13g2_nand3b_1 _11362_ (
    .A_N(addr_i_7_),
    .B(addr_i_5_),
    .C(addr_i_3_),
    .Y(_00981_)
  );
  sg13g2_o21ai_1 _11363_ (
    .A1(_07602_),
    .A2(_03875_),
    .B1(_00981_),
    .Y(_00982_)
  );
  sg13g2_nand2_1 _11364_ (
    .A(addr_i_2_),
    .B(_00982_),
    .Y(_00983_)
  );
  sg13g2_a21oi_1 _11365_ (
    .A1(_00980_),
    .A2(_00983_),
    .B1(addr_i_4_),
    .Y(_00984_)
  );
  sg13g2_nor2_1 _11366_ (
    .A(addr_i_2_),
    .B(_09050_),
    .Y(_00985_)
  );
  sg13g2_o21ai_1 _11367_ (
    .A1(_05236_),
    .A2(_00985_),
    .B1(_00569_),
    .Y(_00986_)
  );
  sg13g2_nor2b_1 _11368_ (
    .A(_00984_),
    .B_N(_00986_),
    .Y(_00987_)
  );
  sg13g2_o21ai_1 _11369_ (
    .A1(addr_i_6_),
    .A2(_00979_),
    .B1(_00987_),
    .Y(_00988_)
  );
  sg13g2_buf_1 _11370_ (
    .A(_05966_),
    .X(_00990_)
  );
  sg13g2_a21oi_1 _11371_ (
    .A1(_00056_),
    .A2(_00368_),
    .B1(addr_i_3_),
    .Y(_00991_)
  );
  sg13g2_a21oi_1 _11372_ (
    .A1(_00990_),
    .A2(_00960_),
    .B1(_00991_),
    .Y(_00992_)
  );
  sg13g2_nor2_1 _11373_ (
    .A(_06386_),
    .B(_01142_),
    .Y(_00993_)
  );
  sg13g2_nand2_1 _11374_ (
    .A(_03435_),
    .B(_04926_),
    .Y(_00994_)
  );
  sg13g2_o21ai_1 _11375_ (
    .A1(_00993_),
    .A2(_03347_),
    .B1(_00994_),
    .Y(_00995_)
  );
  sg13g2_a21oi_1 _11376_ (
    .A1(addr_i_4_),
    .A2(_00995_),
    .B1(_08310_),
    .Y(_00996_)
  );
  sg13g2_o21ai_1 _11377_ (
    .A1(addr_i_2_),
    .A2(_00992_),
    .B1(_00996_),
    .Y(_00997_)
  );
  sg13g2_nor2_1 _11378_ (
    .A(addr_i_3_),
    .B(addr_i_6_),
    .Y(_00998_)
  );
  sg13g2_buf_1 _11379_ (
    .A(_00998_),
    .X(_00999_)
  );
  sg13g2_nand2_1 _11380_ (
    .A(_02602_),
    .B(_00079_),
    .Y(_01001_)
  );
  sg13g2_a21oi_1 _11381_ (
    .A1(_00228_),
    .A2(_02920_),
    .B1(_00059_),
    .Y(_01002_)
  );
  sg13g2_a22oi_1 _11382_ (
    .A1(_00999_),
    .A2(_01001_),
    .B1(_01002_),
    .B2(_09359_),
    .Y(_01003_)
  );
  sg13g2_nand3_1 _11383_ (
    .A(addr_i_2_),
    .B(addr_i_7_),
    .C(addr_i_5_),
    .Y(_01004_)
  );
  sg13g2_nand2_1 _11384_ (
    .A(_00454_),
    .B(_07967_),
    .Y(_01005_)
  );
  sg13g2_o21ai_1 _11385_ (
    .A1(_05745_),
    .A2(_01004_),
    .B1(_01005_),
    .Y(_01006_)
  );
  sg13g2_buf_1 _11386_ (
    .A(_02207_),
    .X(_01007_)
  );
  sg13g2_nand2_1 _11387_ (
    .A(_00637_),
    .B(_04173_),
    .Y(_01008_)
  );
  sg13g2_a21oi_1 _11388_ (
    .A1(_00870_),
    .A2(_01007_),
    .B1(_01008_),
    .Y(_01009_)
  );
  sg13g2_a21oi_1 _11389_ (
    .A1(addr_i_6_),
    .A2(_01006_),
    .B1(_01009_),
    .Y(_01010_)
  );
  sg13g2_o21ai_1 _11390_ (
    .A1(addr_i_7_),
    .A2(_01003_),
    .B1(_01010_),
    .Y(_01012_)
  );
  sg13g2_mux4_1 _11391_ (
    .A0(_00971_),
    .A1(_00988_),
    .A2(_00997_),
    .A3(_01012_),
    .S0(_00113_),
    .S1(addr_i_9_),
    .X(_01013_)
  );
  sg13g2_buf_1 _11392_ (
    .A(_00879_),
    .X(_01014_)
  );
  sg13g2_buf_1 _11393_ (
    .A(_01014_),
    .X(_01015_)
  );
  sg13g2_nor2_1 _11394_ (
    .A(_05910_),
    .B(_08453_),
    .Y(_01016_)
  );
  sg13g2_nor2_1 _11395_ (
    .A(_00687_),
    .B(_00522_),
    .Y(_01017_)
  );
  sg13g2_a22oi_1 _11396_ (
    .A1(_01015_),
    .A2(_00156_),
    .B1(_01016_),
    .B2(_01017_),
    .Y(_01018_)
  );
  sg13g2_buf_1 _11397_ (
    .A(_04151_),
    .X(_01019_)
  );
  sg13g2_nor2_1 _11398_ (
    .A(_06143_),
    .B(_00448_),
    .Y(_01020_)
  );
  sg13g2_nand2_1 _11399_ (
    .A(_01019_),
    .B(_01020_),
    .Y(_01021_)
  );
  sg13g2_o21ai_1 _11400_ (
    .A1(addr_i_5_),
    .A2(_01018_),
    .B1(_01021_),
    .Y(_01023_)
  );
  sg13g2_buf_1 _11401_ (
    .A(_04849_),
    .X(_01024_)
  );
  sg13g2_nor2_1 _11402_ (
    .A(addr_i_3_),
    .B(_00770_),
    .Y(_01025_)
  );
  sg13g2_a21oi_1 _11403_ (
    .A1(addr_i_4_),
    .A2(addr_i_2_),
    .B1(addr_i_6_),
    .Y(_01026_)
  );
  sg13g2_nor3_1 _11404_ (
    .A(_01024_),
    .B(_01025_),
    .C(_01026_),
    .Y(_01027_)
  );
  sg13g2_nand3b_1 _11405_ (
    .A_N(addr_i_6_),
    .B(addr_i_2_),
    .C(addr_i_4_),
    .Y(_01028_)
  );
  sg13g2_buf_1 _11406_ (
    .A(_01028_),
    .X(_01029_)
  );
  sg13g2_nand2_1 _11407_ (
    .A(_00695_),
    .B(_01029_),
    .Y(_01030_)
  );
  sg13g2_buf_1 _11408_ (
    .A(_00721_),
    .X(_01031_)
  );
  sg13g2_a22oi_1 _11409_ (
    .A1(addr_i_3_),
    .A2(_01030_),
    .B1(_01031_),
    .B2(addr_i_5_),
    .Y(_01032_)
  );
  sg13g2_buf_1 _11410_ (
    .A(_07603_),
    .X(_01034_)
  );
  sg13g2_a22oi_1 _11411_ (
    .A1(addr_i_5_),
    .A2(_01027_),
    .B1(_01032_),
    .B2(_01034_),
    .Y(_01035_)
  );
  sg13g2_a21oi_1 _11412_ (
    .A1(_00610_),
    .A2(_01023_),
    .B1(_01035_),
    .Y(_01036_)
  );
  sg13g2_nand2_1 _11413_ (
    .A(_03369_),
    .B(_04860_),
    .Y(_01037_)
  );
  sg13g2_a21oi_1 _11414_ (
    .A1(_00785_),
    .A2(_01037_),
    .B1(addr_i_2_),
    .Y(_01038_)
  );
  sg13g2_a21oi_1 _11415_ (
    .A1(_00594_),
    .A2(_00568_),
    .B1(_01038_),
    .Y(_01039_)
  );
  sg13g2_o21ai_1 _11416_ (
    .A1(_08464_),
    .A2(_08863_),
    .B1(_02250_),
    .Y(_01040_)
  );
  sg13g2_nor2_1 _11417_ (
    .A(_05734_),
    .B(_00019_),
    .Y(_01041_)
  );
  sg13g2_a22oi_1 _11418_ (
    .A1(_04251_),
    .A2(_01040_),
    .B1(_01041_),
    .B2(addr_i_7_),
    .Y(_01042_)
  );
  sg13g2_buf_1 _11419_ (
    .A(_00112_),
    .X(_01043_)
  );
  sg13g2_a22oi_1 _11420_ (
    .A1(addr_i_7_),
    .A2(_01039_),
    .B1(_01042_),
    .B2(_01043_),
    .Y(_01045_)
  );
  sg13g2_nor2_1 _11421_ (
    .A(addr_i_9_),
    .B(_01045_),
    .Y(_01046_)
  );
  sg13g2_nor2_1 _11422_ (
    .A(addr_i_6_),
    .B(_00780_),
    .Y(_01047_)
  );
  sg13g2_nor2_1 _11423_ (
    .A(_02591_),
    .B(_03490_),
    .Y(_01048_)
  );
  sg13g2_buf_1 _11424_ (
    .A(_01048_),
    .X(_01049_)
  );
  sg13g2_nand2_1 _11425_ (
    .A(_05390_),
    .B(_02108_),
    .Y(_01050_)
  );
  sg13g2_a21o_1 _11426_ (
    .A1(_00327_),
    .A2(_01406_),
    .B1(_00637_),
    .X(_01051_)
  );
  sg13g2_a21oi_1 _11427_ (
    .A1(_01050_),
    .A2(_01051_),
    .B1(addr_i_3_),
    .Y(_01052_)
  );
  sg13g2_nor2_1 _11428_ (
    .A(_01049_),
    .B(_01052_),
    .Y(_01053_)
  );
  sg13g2_xor2_1 _11429_ (
    .A(addr_i_2_),
    .B(addr_i_7_),
    .X(_01054_)
  );
  sg13g2_nand2_1 _11430_ (
    .A(_07757_),
    .B(_01054_),
    .Y(_01056_)
  );
  sg13g2_nand2_1 _11431_ (
    .A(addr_i_6_),
    .B(_06851_),
    .Y(_01057_)
  );
  sg13g2_a21oi_1 _11432_ (
    .A1(_01592_),
    .A2(_05910_),
    .B1(addr_i_5_),
    .Y(_01058_)
  );
  sg13g2_a22oi_1 _11433_ (
    .A1(addr_i_7_),
    .A2(_01057_),
    .B1(_01058_),
    .B2(_06419_),
    .Y(_01059_)
  );
  sg13g2_nand2_1 _11434_ (
    .A(_00593_),
    .B(_06530_),
    .Y(_01060_)
  );
  sg13g2_a21oi_1 _11435_ (
    .A1(_00249_),
    .A2(_00549_),
    .B1(_01060_),
    .Y(_01061_)
  );
  sg13g2_a22oi_1 _11436_ (
    .A1(_01056_),
    .A2(_01059_),
    .B1(addr_i_8_),
    .B2(_01061_),
    .Y(_01062_)
  );
  sg13g2_o21ai_1 _11437_ (
    .A1(addr_i_7_),
    .A2(_01053_),
    .B1(_01062_),
    .Y(_01063_)
  );
  sg13g2_nor2_1 _11438_ (
    .A(_03908_),
    .B(_00679_),
    .Y(_01064_)
  );
  sg13g2_buf_1 _11439_ (
    .A(_00678_),
    .X(_01065_)
  );
  sg13g2_buf_1 _11440_ (
    .A(_05324_),
    .X(_01067_)
  );
  sg13g2_a21oi_1 _11441_ (
    .A1(_06862_),
    .A2(_01065_),
    .B1(_01067_),
    .Y(_01068_)
  );
  sg13g2_o21ai_1 _11442_ (
    .A1(_01064_),
    .A2(_01068_),
    .B1(addr_i_6_),
    .Y(_01069_)
  );
  sg13g2_buf_1 _11443_ (
    .A(_08376_),
    .X(_01070_)
  );
  sg13g2_nand3_1 _11444_ (
    .A(_01070_),
    .B(_00376_),
    .C(_00320_),
    .Y(_01071_)
  );
  sg13g2_a21oi_1 _11445_ (
    .A1(_01768_),
    .A2(_02920_),
    .B1(addr_i_3_),
    .Y(_01072_)
  );
  sg13g2_nand2_1 _11446_ (
    .A(addr_i_3_),
    .B(_03106_),
    .Y(_01073_)
  );
  sg13g2_a21oi_1 _11447_ (
    .A1(_00878_),
    .A2(_01073_),
    .B1(addr_i_5_),
    .Y(_01074_)
  );
  sg13g2_o21ai_1 _11448_ (
    .A1(_01072_),
    .A2(_01074_),
    .B1(addr_i_7_),
    .Y(_01075_)
  );
  sg13g2_nand4_1 _11449_ (
    .A(addr_i_8_),
    .B(_01069_),
    .C(_01071_),
    .D(_01075_),
    .Y(_01076_)
  );
  sg13g2_a221oi_1 _11450_ (
    .A1(_01047_),
    .A2(_00503_),
    .B1(_01063_),
    .B2(_01076_),
    .C1(_01351_),
    .Y(_01078_)
  );
  sg13g2_a22oi_1 _11451_ (
    .A1(_01036_),
    .A2(_01046_),
    .B1(addr_i_10_),
    .B2(_01078_),
    .Y(_01079_)
  );
  sg13g2_a22oi_1 _11452_ (
    .A1(addr_i_10_),
    .A2(_01013_),
    .B1(_01079_),
    .B2(addr_i_11_),
    .Y(_01080_)
  );
  sg13g2_a22oi_1 _11453_ (
    .A1(_00891_),
    .A2(_00958_),
    .B1(addr_i_12_),
    .B2(_01080_),
    .Y(_01081_)
  );
  sg13g2_or2_1 _11454_ (
    .A(_00814_),
    .B(_01081_),
    .X(data_o_11_)
  );
  sg13g2_buf_1 _11455_ (
    .A(_00860_),
    .X(_01082_)
  );
  sg13g2_nand3_1 _11456_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .C(addr_i_5_),
    .Y(_01083_)
  );
  sg13g2_buf_1 _11457_ (
    .A(_01083_),
    .X(_01084_)
  );
  sg13g2_nand2_1 _11458_ (
    .A(_00878_),
    .B(_01084_),
    .Y(_01085_)
  );
  sg13g2_buf_1 _11459_ (
    .A(_03128_),
    .X(_01086_)
  );
  sg13g2_o21ai_1 _11460_ (
    .A1(addr_i_3_),
    .A2(_01086_),
    .B1(_00261_),
    .Y(_01088_)
  );
  sg13g2_nand3_1 _11461_ (
    .A(_00115_),
    .B(addr_i_6_),
    .C(_06032_),
    .Y(_01089_)
  );
  sg13g2_a21oi_1 _11462_ (
    .A1(_01088_),
    .A2(_01089_),
    .B1(addr_i_5_),
    .Y(_01090_)
  );
  sg13g2_nor2_1 _11463_ (
    .A(_04418_),
    .B(_00406_),
    .Y(_01091_)
  );
  sg13g2_a22oi_1 _11464_ (
    .A1(addr_i_3_),
    .A2(_01085_),
    .B1(_01090_),
    .B2(_01091_),
    .Y(_01092_)
  );
  sg13g2_nor2_1 _11465_ (
    .A(addr_i_3_),
    .B(_01965_),
    .Y(_01093_)
  );
  sg13g2_nor2_1 _11466_ (
    .A(addr_i_2_),
    .B(_06530_),
    .Y(_01094_)
  );
  sg13g2_buf_1 _11467_ (
    .A(_00343_),
    .X(_01095_)
  );
  sg13g2_o21ai_1 _11468_ (
    .A1(_01093_),
    .A2(_01094_),
    .B1(_01095_),
    .Y(_01096_)
  );
  sg13g2_nand2_1 _11469_ (
    .A(_03765_),
    .B(_00078_),
    .Y(_01097_)
  );
  sg13g2_buf_1 _11470_ (
    .A(_00780_),
    .X(_01099_)
  );
  sg13g2_a22oi_1 _11471_ (
    .A1(_00999_),
    .A2(_01097_),
    .B1(_01099_),
    .B2(_00743_),
    .Y(_01100_)
  );
  sg13g2_nand3b_1 _11472_ (
    .A_N(_00369_),
    .B(_01096_),
    .C(_01100_),
    .Y(_01101_)
  );
  sg13g2_o21ai_1 _11473_ (
    .A1(_01082_),
    .A2(_01092_),
    .B1(_01101_),
    .Y(_01102_)
  );
  sg13g2_buf_1 _11474_ (
    .A(_03875_),
    .X(_01103_)
  );
  sg13g2_buf_1 _11475_ (
    .A(_00024_),
    .X(_01104_)
  );
  sg13g2_a21oi_1 _11476_ (
    .A1(_00659_),
    .A2(_01103_),
    .B1(_01104_),
    .Y(_01105_)
  );
  sg13g2_nor2_1 _11477_ (
    .A(addr_i_4_),
    .B(_00451_),
    .Y(_01106_)
  );
  sg13g2_buf_1 _11478_ (
    .A(_01106_),
    .X(_01107_)
  );
  sg13g2_o21ai_1 _11479_ (
    .A1(_00244_),
    .A2(_01107_),
    .B1(addr_i_3_),
    .Y(_01108_)
  );
  sg13g2_a21oi_1 _11480_ (
    .A1(_06508_),
    .A2(_01108_),
    .B1(addr_i_6_),
    .Y(_01110_)
  );
  sg13g2_a22oi_1 _11481_ (
    .A1(_00073_),
    .A2(_00329_),
    .B1(_01105_),
    .B2(_01110_),
    .Y(_01111_)
  );
  sg13g2_buf_1 _11482_ (
    .A(_00934_),
    .X(_01112_)
  );
  sg13g2_buf_1 _11483_ (
    .A(_07933_),
    .X(_01113_)
  );
  sg13g2_buf_1 _11484_ (
    .A(_01113_),
    .X(_01114_)
  );
  sg13g2_o21ai_1 _11485_ (
    .A1(_01112_),
    .A2(_06264_),
    .B1(_01114_),
    .Y(_01115_)
  );
  sg13g2_a21oi_1 _11486_ (
    .A1(_00907_),
    .A2(_01115_),
    .B1(addr_i_3_),
    .Y(_01116_)
  );
  sg13g2_nor3_1 _11487_ (
    .A(_07547_),
    .B(_00409_),
    .C(_00626_),
    .Y(_01117_)
  );
  sg13g2_buf_1 _11488_ (
    .A(_07934_),
    .X(_01118_)
  );
  sg13g2_buf_1 _11489_ (
    .A(_01118_),
    .X(_01119_)
  );
  sg13g2_o21ai_1 _11490_ (
    .A1(_01116_),
    .A2(_01117_),
    .B1(_01119_),
    .Y(_01121_)
  );
  sg13g2_o21ai_1 _11491_ (
    .A1(_03238_),
    .A2(_01111_),
    .B1(_01121_),
    .Y(_01122_)
  );
  sg13g2_or2_1 _11492_ (
    .A(_01102_),
    .B(_01122_),
    .X(_01123_)
  );
  sg13g2_nor2_1 _11493_ (
    .A(addr_i_10_),
    .B(_00397_),
    .Y(_01124_)
  );
  sg13g2_buf_1 _11494_ (
    .A(_05036_),
    .X(_01125_)
  );
  sg13g2_nand2_1 _11495_ (
    .A(_04296_),
    .B(_01125_),
    .Y(_01126_)
  );
  sg13g2_nor2_1 _11496_ (
    .A(addr_i_2_),
    .B(_00678_),
    .Y(_01127_)
  );
  sg13g2_nor2_1 _11497_ (
    .A(_06298_),
    .B(_01127_),
    .Y(_01128_)
  );
  sg13g2_nor2_1 _11498_ (
    .A(addr_i_4_),
    .B(_01128_),
    .Y(_01129_)
  );
  sg13g2_a22oi_1 _11499_ (
    .A1(addr_i_4_),
    .A2(_01126_),
    .B1(_01129_),
    .B2(_06740_),
    .Y(_01130_)
  );
  sg13g2_nand2_1 _11500_ (
    .A(_00377_),
    .B(_00818_),
    .Y(_01132_)
  );
  sg13g2_o21ai_1 _11501_ (
    .A1(addr_i_3_),
    .A2(_01130_),
    .B1(_01132_),
    .Y(_01133_)
  );
  sg13g2_nand2_1 _11502_ (
    .A(_03953_),
    .B(_00981_),
    .Y(_01134_)
  );
  sg13g2_a21o_1 _11503_ (
    .A1(addr_i_4_),
    .A2(_01134_),
    .B1(_04506_),
    .X(_01135_)
  );
  sg13g2_a221oi_1 _11504_ (
    .A1(addr_i_6_),
    .A2(_01133_),
    .B1(_01135_),
    .B2(addr_i_2_),
    .C1(addr_i_8_),
    .Y(_01136_)
  );
  sg13g2_nand2_1 _11505_ (
    .A(_09486_),
    .B(_08598_),
    .Y(_01137_)
  );
  sg13g2_nor2_1 _11506_ (
    .A(_00070_),
    .B(_02755_),
    .Y(_01138_)
  );
  sg13g2_nor2_1 _11507_ (
    .A(_00150_),
    .B(_06927_),
    .Y(_01139_)
  );
  sg13g2_o21ai_1 _11508_ (
    .A1(_01138_),
    .A2(_01139_),
    .B1(_00388_),
    .Y(_01140_)
  );
  sg13g2_a21oi_1 _11509_ (
    .A1(_01137_),
    .A2(_01140_),
    .B1(addr_i_3_),
    .Y(_01141_)
  );
  sg13g2_a21oi_1 _11510_ (
    .A1(addr_i_5_),
    .A2(_09492_),
    .B1(_00531_),
    .Y(_01143_)
  );
  sg13g2_buf_1 _11511_ (
    .A(_01197_),
    .X(_01144_)
  );
  sg13g2_a21oi_1 _11512_ (
    .A1(_00051_),
    .A2(_01144_),
    .B1(addr_i_4_),
    .Y(_01145_)
  );
  sg13g2_o21ai_1 _11513_ (
    .A1(_01143_),
    .A2(_01145_),
    .B1(addr_i_2_),
    .Y(_01146_)
  );
  sg13g2_nand2_1 _11514_ (
    .A(addr_i_6_),
    .B(_00069_),
    .Y(_01147_)
  );
  sg13g2_or2_1 _11515_ (
    .A(_05490_),
    .B(_01147_),
    .X(_01148_)
  );
  sg13g2_nand3_1 _11516_ (
    .A(addr_i_8_),
    .B(_01146_),
    .C(_01148_),
    .Y(_01149_)
  );
  sg13g2_o21ai_1 _11517_ (
    .A1(_01141_),
    .A2(_01149_),
    .B1(_00773_),
    .Y(_01150_)
  );
  sg13g2_buf_1 _11518_ (
    .A(_01559_),
    .X(_01151_)
  );
  sg13g2_nand2_1 _11519_ (
    .A(addr_i_5_),
    .B(_01669_),
    .Y(_01152_)
  );
  sg13g2_nand2_1 _11520_ (
    .A(_04384_),
    .B(_01152_),
    .Y(_01154_)
  );
  sg13g2_buf_1 _11521_ (
    .A(_00316_),
    .X(_01155_)
  );
  sg13g2_o21ai_1 _11522_ (
    .A1(_05811_),
    .A2(_01086_),
    .B1(addr_i_2_),
    .Y(_01156_)
  );
  sg13g2_a21oi_1 _11523_ (
    .A1(_01155_),
    .A2(_01156_),
    .B1(addr_i_5_),
    .Y(_01157_)
  );
  sg13g2_a22oi_1 _11524_ (
    .A1(addr_i_4_),
    .A2(_01154_),
    .B1(_01157_),
    .B2(addr_i_3_),
    .Y(_01158_)
  );
  sg13g2_buf_1 _11525_ (
    .A(_01680_),
    .X(_01159_)
  );
  sg13g2_buf_1 _11526_ (
    .A(_06851_),
    .X(_01160_)
  );
  sg13g2_o21ai_1 _11527_ (
    .A1(_01159_),
    .A2(_01160_),
    .B1(_00077_),
    .Y(_01161_)
  );
  sg13g2_o21ai_1 _11528_ (
    .A1(_00688_),
    .A2(_00448_),
    .B1(_00704_),
    .Y(_01162_)
  );
  sg13g2_nand2_1 _11529_ (
    .A(addr_i_3_),
    .B(_00655_),
    .Y(_01163_)
  );
  sg13g2_a221oi_1 _11530_ (
    .A1(addr_i_5_),
    .A2(_01161_),
    .B1(_01162_),
    .B2(addr_i_7_),
    .C1(_01163_),
    .Y(_01165_)
  );
  sg13g2_nor3_1 _11531_ (
    .A(_01151_),
    .B(_01158_),
    .C(_01165_),
    .Y(_01166_)
  );
  sg13g2_nand2_1 _11532_ (
    .A(_02920_),
    .B(_00368_),
    .Y(_01167_)
  );
  sg13g2_nand2_1 _11533_ (
    .A(_05390_),
    .B(_00000_),
    .Y(_01168_)
  );
  sg13g2_buf_1 _11534_ (
    .A(_01067_),
    .X(_01169_)
  );
  sg13g2_a21oi_1 _11535_ (
    .A1(_00567_),
    .A2(_01168_),
    .B1(_01169_),
    .Y(_01170_)
  );
  sg13g2_a22oi_1 _11536_ (
    .A1(_00116_),
    .A2(_01167_),
    .B1(_01170_),
    .B2(_01049_),
    .Y(_01171_)
  );
  sg13g2_nand4_1 _11537_ (
    .A(_00703_),
    .B(_01047_),
    .C(_00105_),
    .D(_00344_),
    .Y(_01172_)
  );
  sg13g2_o21ai_1 _11538_ (
    .A1(_01082_),
    .A2(_01171_),
    .B1(_01172_),
    .Y(_01173_)
  );
  sg13g2_nor2_1 _11539_ (
    .A(_03731_),
    .B(addr_i_9_),
    .Y(_01174_)
  );
  sg13g2_buf_1 _11540_ (
    .A(_01174_),
    .X(_01176_)
  );
  sg13g2_o21ai_1 _11541_ (
    .A1(_01166_),
    .A2(_01173_),
    .B1(_01176_),
    .Y(_01177_)
  );
  sg13g2_o21ai_1 _11542_ (
    .A1(_01136_),
    .A2(_01150_),
    .B1(_01177_),
    .Y(_01178_)
  );
  sg13g2_buf_1 _11543_ (
    .A(_00038_),
    .X(_01179_)
  );
  sg13g2_nand2_1 _11544_ (
    .A(_00428_),
    .B(_00375_),
    .Y(_01180_)
  );
  sg13g2_o21ai_1 _11545_ (
    .A1(_01179_),
    .A2(_01180_),
    .B1(addr_i_8_),
    .Y(_01181_)
  );
  sg13g2_nand2_1 _11546_ (
    .A(addr_i_3_),
    .B(_04086_),
    .Y(_01182_)
  );
  sg13g2_nand2_1 _11547_ (
    .A(_00731_),
    .B(_01182_),
    .Y(_01183_)
  );
  sg13g2_nor2_1 _11548_ (
    .A(addr_i_3_),
    .B(_01179_),
    .Y(_01184_)
  );
  sg13g2_a21oi_1 _11549_ (
    .A1(addr_i_4_),
    .A2(_01183_),
    .B1(_01184_),
    .Y(_01185_)
  );
  sg13g2_a21oi_1 _11550_ (
    .A1(_02799_),
    .A2(_02634_),
    .B1(_00059_),
    .Y(_01187_)
  );
  sg13g2_o21ai_1 _11551_ (
    .A1(_01041_),
    .A2(_01187_),
    .B1(_00529_),
    .Y(_01188_)
  );
  sg13g2_o21ai_1 _11552_ (
    .A1(_00390_),
    .A2(_01185_),
    .B1(_01188_),
    .Y(_01189_)
  );
  sg13g2_o21ai_1 _11553_ (
    .A1(_01181_),
    .A2(_01189_),
    .B1(_05203_),
    .Y(_01190_)
  );
  sg13g2_buf_1 _11554_ (
    .A(_00165_),
    .X(_01191_)
  );
  sg13g2_nor2_1 _11555_ (
    .A(addr_i_3_),
    .B(_07602_),
    .Y(_01192_)
  );
  sg13g2_nor2_1 _11556_ (
    .A(_01191_),
    .B(_01192_),
    .Y(_01193_)
  );
  sg13g2_buf_1 _11557_ (
    .A(_04782_),
    .X(_01194_)
  );
  sg13g2_o21ai_1 _11558_ (
    .A1(_06795_),
    .A2(_01194_),
    .B1(addr_i_3_),
    .Y(_01195_)
  );
  sg13g2_a21o_1 _11559_ (
    .A1(_09149_),
    .A2(_01195_),
    .B1(_08399_),
    .X(_01196_)
  );
  sg13g2_o21ai_1 _11560_ (
    .A1(_06873_),
    .A2(_01193_),
    .B1(_01196_),
    .Y(_01198_)
  );
  sg13g2_nand2_1 _11561_ (
    .A(_07381_),
    .B(_04173_),
    .Y(_01199_)
  );
  sg13g2_a21oi_1 _11562_ (
    .A1(_01199_),
    .A2(_00077_),
    .B1(addr_i_3_),
    .Y(_01200_)
  );
  sg13g2_a21oi_1 _11563_ (
    .A1(_00529_),
    .A2(_00818_),
    .B1(_01200_),
    .Y(_01201_)
  );
  sg13g2_nor2_1 _11564_ (
    .A(_03908_),
    .B(_02722_),
    .Y(_01202_)
  );
  sg13g2_buf_1 _11565_ (
    .A(_04395_),
    .X(_01203_)
  );
  sg13g2_a22oi_1 _11566_ (
    .A1(_01203_),
    .A2(_00747_),
    .B1(_00157_),
    .B2(addr_i_6_),
    .Y(_01204_)
  );
  sg13g2_a22oi_1 _11567_ (
    .A1(_00029_),
    .A2(_01202_),
    .B1(_01204_),
    .B2(addr_i_8_),
    .Y(_01205_)
  );
  sg13g2_o21ai_1 _11568_ (
    .A1(addr_i_5_),
    .A2(_01201_),
    .B1(_01205_),
    .Y(_01206_)
  );
  sg13g2_a21oi_1 _11569_ (
    .A1(addr_i_6_),
    .A2(_01198_),
    .B1(_01206_),
    .Y(_01207_)
  );
  sg13g2_o21ai_1 _11570_ (
    .A1(_01190_),
    .A2(_01207_),
    .B1(_00312_),
    .Y(_01209_)
  );
  sg13g2_a22oi_1 _11571_ (
    .A1(_01123_),
    .A2(_01124_),
    .B1(_01178_),
    .B2(_01209_),
    .Y(_01210_)
  );
  sg13g2_buf_1 _11572_ (
    .A(_03073_),
    .X(_01211_)
  );
  sg13g2_buf_1 _11573_ (
    .A(_00246_),
    .X(_01212_)
  );
  sg13g2_nand2_1 _11574_ (
    .A(_01212_),
    .B(_00764_),
    .Y(_01213_)
  );
  sg13g2_a22oi_1 _11575_ (
    .A1(_00305_),
    .A2(_01213_),
    .B1(_00436_),
    .B2(addr_i_3_),
    .Y(_01214_)
  );
  sg13g2_buf_1 _11576_ (
    .A(_07956_),
    .X(_01215_)
  );
  sg13g2_buf_1 _11577_ (
    .A(_01215_),
    .X(_01216_)
  );
  sg13g2_a22oi_1 _11578_ (
    .A1(addr_i_5_),
    .A2(_00578_),
    .B1(_01216_),
    .B2(_01024_),
    .Y(_01217_)
  );
  sg13g2_a21oi_1 _11579_ (
    .A1(_03964_),
    .A2(_01217_),
    .B1(_00191_),
    .Y(_01218_)
  );
  sg13g2_nor2_1 _11580_ (
    .A(_01214_),
    .B(_01218_),
    .Y(_01220_)
  );
  sg13g2_nand2_1 _11581_ (
    .A(_00176_),
    .B(_00000_),
    .Y(_01221_)
  );
  sg13g2_buf_1 _11582_ (
    .A(_01221_),
    .X(_01222_)
  );
  sg13g2_nand2_1 _11583_ (
    .A(_00516_),
    .B(_01222_),
    .Y(_01223_)
  );
  sg13g2_buf_1 _11584_ (
    .A(_00863_),
    .X(_01224_)
  );
  sg13g2_a21oi_1 _11585_ (
    .A1(_03391_),
    .A2(_01224_),
    .B1(addr_i_7_),
    .Y(_01225_)
  );
  sg13g2_a22oi_1 _11586_ (
    .A1(addr_i_3_),
    .A2(_01223_),
    .B1(_01225_),
    .B2(addr_i_2_),
    .Y(_01226_)
  );
  sg13g2_buf_1 _11587_ (
    .A(_07458_),
    .X(_01227_)
  );
  sg13g2_xnor2_1 _11588_ (
    .A(addr_i_7_),
    .B(addr_i_5_),
    .Y(_01228_)
  );
  sg13g2_nor2_1 _11589_ (
    .A(addr_i_7_),
    .B(_04793_),
    .Y(_01229_)
  );
  sg13g2_buf_1 _11590_ (
    .A(_01229_),
    .X(_01231_)
  );
  sg13g2_buf_1 _11591_ (
    .A(_00897_),
    .X(_01232_)
  );
  sg13g2_o21ai_1 _11592_ (
    .A1(_01231_),
    .A2(_01232_),
    .B1(_08752_),
    .Y(_01233_)
  );
  sg13g2_nand2_1 _11593_ (
    .A(addr_i_3_),
    .B(_04284_),
    .Y(_01234_)
  );
  sg13g2_a21oi_1 _11594_ (
    .A1(_01233_),
    .A2(_01234_),
    .B1(addr_i_4_),
    .Y(_01235_)
  );
  sg13g2_a22oi_1 _11595_ (
    .A1(_01227_),
    .A2(_01228_),
    .B1(_01235_),
    .B2(_00123_),
    .Y(_01236_)
  );
  sg13g2_nor3_1 _11596_ (
    .A(_03259_),
    .B(_01226_),
    .C(_01236_),
    .Y(_01237_)
  );
  sg13g2_a21oi_1 _11597_ (
    .A1(_00114_),
    .A2(_01220_),
    .B1(_01237_),
    .Y(_01238_)
  );
  sg13g2_nor2_1 _11598_ (
    .A(_01211_),
    .B(_01238_),
    .Y(_01239_)
  );
  sg13g2_buf_1 _11599_ (
    .A(_07503_),
    .X(_01240_)
  );
  sg13g2_a21oi_1 _11600_ (
    .A1(_00022_),
    .A2(_01227_),
    .B1(_01240_),
    .Y(_01242_)
  );
  sg13g2_nor2b_1 _11601_ (
    .A(addr_i_3_),
    .B_N(addr_i_5_),
    .Y(_01243_)
  );
  sg13g2_buf_1 _11602_ (
    .A(_01243_),
    .X(_01244_)
  );
  sg13g2_nand2_1 _11603_ (
    .A(_08564_),
    .B(_01244_),
    .Y(_01245_)
  );
  sg13g2_nor2_1 _11604_ (
    .A(_08741_),
    .B(_00770_),
    .Y(_01246_)
  );
  sg13g2_o21ai_1 _11605_ (
    .A1(_00031_),
    .A2(_01246_),
    .B1(_06154_),
    .Y(_01247_)
  );
  sg13g2_a21o_1 _11606_ (
    .A1(_01245_),
    .A2(_01247_),
    .B1(addr_i_6_),
    .X(_01248_)
  );
  sg13g2_o21ai_1 _11607_ (
    .A1(_00123_),
    .A2(_01242_),
    .B1(_01248_),
    .Y(_01249_)
  );
  sg13g2_a22oi_1 _11608_ (
    .A1(_00485_),
    .A2(_00414_),
    .B1(addr_i_5_),
    .B2(addr_i_4_),
    .Y(_01250_)
  );
  sg13g2_a21oi_1 _11609_ (
    .A1(addr_i_4_),
    .A2(_00941_),
    .B1(_01250_),
    .Y(_01251_)
  );
  sg13g2_o21ai_1 _11610_ (
    .A1(_01034_),
    .A2(_01251_),
    .B1(addr_i_9_),
    .Y(_01253_)
  );
  sg13g2_o21ai_1 _11611_ (
    .A1(addr_i_4_),
    .A2(_01066_),
    .B1(_00327_),
    .Y(_01254_)
  );
  sg13g2_nor2_1 _11612_ (
    .A(_06364_),
    .B(_05524_),
    .Y(_01255_)
  );
  sg13g2_o21ai_1 _11613_ (
    .A1(addr_i_5_),
    .A2(_01255_),
    .B1(_00704_),
    .Y(_01256_)
  );
  sg13g2_buf_1 _11614_ (
    .A(_00327_),
    .X(_01257_)
  );
  sg13g2_o21ai_1 _11615_ (
    .A1(addr_i_6_),
    .A2(_00269_),
    .B1(addr_i_4_),
    .Y(_01258_)
  );
  sg13g2_a21oi_1 _11616_ (
    .A1(_01257_),
    .A2(_01258_),
    .B1(addr_i_7_),
    .Y(_01259_)
  );
  sg13g2_a221oi_1 _11617_ (
    .A1(addr_i_5_),
    .A2(_01254_),
    .B1(_01256_),
    .B2(addr_i_7_),
    .C1(_01259_),
    .Y(_01260_)
  );
  sg13g2_inv_1 _11618_ (
    .A(_01260_),
    .Y(_01261_)
  );
  sg13g2_buf_1 _11619_ (
    .A(_00297_),
    .X(_01262_)
  );
  sg13g2_nand2_1 _11620_ (
    .A(_06840_),
    .B(_03709_),
    .Y(_01264_)
  );
  sg13g2_nand2_1 _11621_ (
    .A(_00676_),
    .B(_03194_),
    .Y(_01265_)
  );
  sg13g2_nand2_1 _11622_ (
    .A(_00701_),
    .B(_01265_),
    .Y(_01266_)
  );
  sg13g2_nand2_1 _11623_ (
    .A(_02152_),
    .B(_00252_),
    .Y(_01267_)
  );
  sg13g2_nand2_1 _11624_ (
    .A(addr_i_5_),
    .B(_00768_),
    .Y(_01268_)
  );
  sg13g2_a21oi_1 _11625_ (
    .A1(_01267_),
    .A2(_01268_),
    .B1(addr_i_7_),
    .Y(_01269_)
  );
  sg13g2_a22oi_1 _11626_ (
    .A1(_01262_),
    .A2(_01264_),
    .B1(_01266_),
    .B2(_01269_),
    .Y(_01270_)
  );
  sg13g2_a22oi_1 _11627_ (
    .A1(addr_i_3_),
    .A2(_01261_),
    .B1(_01270_),
    .B2(_03259_),
    .Y(_01271_)
  );
  sg13g2_a22oi_1 _11628_ (
    .A1(_00277_),
    .A2(_01249_),
    .B1(_01253_),
    .B2(_01271_),
    .Y(_01272_)
  );
  sg13g2_buf_1 _11629_ (
    .A(_07469_),
    .X(_01273_)
  );
  sg13g2_nand2_1 _11630_ (
    .A(_01113_),
    .B(_01273_),
    .Y(_01275_)
  );
  sg13g2_buf_1 _11631_ (
    .A(_04749_),
    .X(_01276_)
  );
  sg13g2_buf_1 _11632_ (
    .A(_01276_),
    .X(_01277_)
  );
  sg13g2_nor3_1 _11633_ (
    .A(addr_i_3_),
    .B(_01277_),
    .C(_00559_),
    .Y(_01278_)
  );
  sg13g2_buf_1 _11634_ (
    .A(_00445_),
    .X(_01279_)
  );
  sg13g2_a22oi_1 _11635_ (
    .A1(addr_i_3_),
    .A2(_01275_),
    .B1(_01278_),
    .B2(_01279_),
    .Y(_01280_)
  );
  sg13g2_nor2_1 _11636_ (
    .A(_05845_),
    .B(_03709_),
    .Y(_01281_)
  );
  sg13g2_buf_1 _11637_ (
    .A(_00269_),
    .X(_01282_)
  );
  sg13g2_o21ai_1 _11638_ (
    .A1(_06806_),
    .A2(_01281_),
    .B1(_01282_),
    .Y(_01283_)
  );
  sg13g2_nand2b_1 _11639_ (
    .A_N(_01280_),
    .B(_01283_),
    .Y(_01284_)
  );
  sg13g2_nor2_1 _11640_ (
    .A(_00650_),
    .B(_03743_),
    .Y(_01286_)
  );
  sg13g2_nand3_1 _11641_ (
    .A(addr_i_3_),
    .B(_00024_),
    .C(_05457_),
    .Y(_01287_)
  );
  sg13g2_a21oi_1 _11642_ (
    .A1(_00228_),
    .A2(_01287_),
    .B1(_06717_),
    .Y(_01288_)
  );
  sg13g2_o21ai_1 _11643_ (
    .A1(_01286_),
    .A2(_01288_),
    .B1(addr_i_7_),
    .Y(_01289_)
  );
  sg13g2_buf_1 _11644_ (
    .A(_01768_),
    .X(_01290_)
  );
  sg13g2_nand2_1 _11645_ (
    .A(_01104_),
    .B(_01290_),
    .Y(_01291_)
  );
  sg13g2_nor2_1 _11646_ (
    .A(_07381_),
    .B(_00198_),
    .Y(_01292_)
  );
  sg13g2_o21ai_1 _11647_ (
    .A1(_01292_),
    .A2(_00257_),
    .B1(addr_i_3_),
    .Y(_01293_)
  );
  sg13g2_nor2_1 _11648_ (
    .A(_00117_),
    .B(_01680_),
    .Y(_01294_)
  );
  sg13g2_nor2_1 _11649_ (
    .A(_00914_),
    .B(_02426_),
    .Y(_01295_)
  );
  sg13g2_a21oi_1 _11650_ (
    .A1(_00322_),
    .A2(_01294_),
    .B1(_01295_),
    .Y(_01297_)
  );
  sg13g2_a21oi_1 _11651_ (
    .A1(_01293_),
    .A2(_01297_),
    .B1(addr_i_4_),
    .Y(_01298_)
  );
  sg13g2_a21oi_1 _11652_ (
    .A1(_00234_),
    .A2(_01291_),
    .B1(_01298_),
    .Y(_01299_)
  );
  sg13g2_a21oi_1 _11653_ (
    .A1(_01289_),
    .A2(_01299_),
    .B1(addr_i_8_),
    .Y(_01300_)
  );
  sg13g2_buf_1 _11654_ (
    .A(_00915_),
    .X(_01301_)
  );
  sg13g2_buf_1 _11655_ (
    .A(_03665_),
    .X(_01302_)
  );
  sg13g2_a21oi_1 _11656_ (
    .A1(_01301_),
    .A2(_01302_),
    .B1(_00073_),
    .Y(_01303_)
  );
  sg13g2_nor2_1 _11657_ (
    .A(addr_i_5_),
    .B(_00375_),
    .Y(_01304_)
  );
  sg13g2_o21ai_1 _11658_ (
    .A1(addr_i_4_),
    .A2(addr_i_2_),
    .B1(addr_i_5_),
    .Y(_01305_)
  );
  sg13g2_nor2_1 _11659_ (
    .A(addr_i_6_),
    .B(_01305_),
    .Y(_01306_)
  );
  sg13g2_buf_1 _11660_ (
    .A(_00260_),
    .X(_01308_)
  );
  sg13g2_nand2_1 _11661_ (
    .A(_00030_),
    .B(_02722_),
    .Y(_01309_)
  );
  sg13g2_buf_1 _11662_ (
    .A(_00713_),
    .X(_01310_)
  );
  sg13g2_o21ai_1 _11663_ (
    .A1(_01308_),
    .A2(_01309_),
    .B1(_01310_),
    .Y(_01311_)
  );
  sg13g2_a22oi_1 _11664_ (
    .A1(addr_i_6_),
    .A2(_01304_),
    .B1(_01306_),
    .B2(_01311_),
    .Y(_01312_)
  );
  sg13g2_o21ai_1 _11665_ (
    .A1(addr_i_2_),
    .A2(_01303_),
    .B1(_01312_),
    .Y(_01313_)
  );
  sg13g2_nand2_1 _11666_ (
    .A(_00396_),
    .B(_01313_),
    .Y(_01314_)
  );
  sg13g2_a22oi_1 _11667_ (
    .A1(_01119_),
    .A2(_01284_),
    .B1(_01300_),
    .B2(_01314_),
    .Y(_01315_)
  );
  sg13g2_nor3_1 _11668_ (
    .A(addr_i_10_),
    .B(_01272_),
    .C(_01315_),
    .Y(_01316_)
  );
  sg13g2_nand2_1 _11669_ (
    .A(_00223_),
    .B(_09138_),
    .Y(_01317_)
  );
  sg13g2_buf_1 _11670_ (
    .A(_04173_),
    .X(_01319_)
  );
  sg13g2_buf_1 _11671_ (
    .A(_01319_),
    .X(_01320_)
  );
  sg13g2_o21ai_1 _11672_ (
    .A1(_01320_),
    .A2(_00257_),
    .B1(addr_i_3_),
    .Y(_01321_)
  );
  sg13g2_a21oi_1 _11673_ (
    .A1(_01317_),
    .A2(_01321_),
    .B1(addr_i_4_),
    .Y(_01322_)
  );
  sg13g2_nor2_1 _11674_ (
    .A(_00703_),
    .B(_00390_),
    .Y(_01323_)
  );
  sg13g2_buf_1 _11675_ (
    .A(_08708_),
    .X(_01324_)
  );
  sg13g2_o21ai_1 _11676_ (
    .A1(_01322_),
    .A2(_01323_),
    .B1(_01324_),
    .Y(_01325_)
  );
  sg13g2_nand2_1 _11677_ (
    .A(addr_i_6_),
    .B(_00246_),
    .Y(_01326_)
  );
  sg13g2_a21oi_1 _11678_ (
    .A1(addr_i_5_),
    .A2(_01326_),
    .B1(_01015_),
    .Y(_01327_)
  );
  sg13g2_nor2_1 _11679_ (
    .A(addr_i_3_),
    .B(_01327_),
    .Y(_01328_)
  );
  sg13g2_nor2_1 _11680_ (
    .A(_08100_),
    .B(_00977_),
    .Y(_01330_)
  );
  sg13g2_nand2_1 _11681_ (
    .A(_00269_),
    .B(_01867_),
    .Y(_01331_)
  );
  sg13g2_o21ai_1 _11682_ (
    .A1(_00531_),
    .A2(_01330_),
    .B1(_01331_),
    .Y(_01332_)
  );
  sg13g2_or2_1 _11683_ (
    .A(_01328_),
    .B(_01332_),
    .X(_01333_)
  );
  sg13g2_nor2_1 _11684_ (
    .A(_01324_),
    .B(_01180_),
    .Y(_01334_)
  );
  sg13g2_a22oi_1 _11685_ (
    .A1(addr_i_4_),
    .A2(_01333_),
    .B1(_01334_),
    .B2(_00114_),
    .Y(_01335_)
  );
  sg13g2_buf_1 _11686_ (
    .A(_00322_),
    .X(_01336_)
  );
  sg13g2_nand3b_1 _11687_ (
    .A_N(addr_i_5_),
    .B(addr_i_6_),
    .C(addr_i_7_),
    .Y(_01337_)
  );
  sg13g2_nand2_1 _11688_ (
    .A(_00679_),
    .B(_01337_),
    .Y(_01338_)
  );
  sg13g2_buf_1 _11689_ (
    .A(_02196_),
    .X(_01339_)
  );
  sg13g2_a21oi_1 _11690_ (
    .A1(_03964_),
    .A2(_00051_),
    .B1(_01339_),
    .Y(_01341_)
  );
  sg13g2_a21oi_1 _11691_ (
    .A1(_00239_),
    .A2(_01338_),
    .B1(_01341_),
    .Y(_01342_)
  );
  sg13g2_buf_1 _11692_ (
    .A(_00620_),
    .X(_01343_)
  );
  sg13g2_a21oi_1 _11693_ (
    .A1(_06784_),
    .A2(_01343_),
    .B1(addr_i_3_),
    .Y(_01344_)
  );
  sg13g2_a22oi_1 _11694_ (
    .A1(_01282_),
    .A2(_00529_),
    .B1(_01344_),
    .B2(addr_i_4_),
    .Y(_01345_)
  );
  sg13g2_a21oi_1 _11695_ (
    .A1(addr_i_4_),
    .A2(_01342_),
    .B1(_01345_),
    .Y(_01346_)
  );
  sg13g2_a22oi_1 _11696_ (
    .A1(_01336_),
    .A2(_00898_),
    .B1(_01346_),
    .B2(addr_i_8_),
    .Y(_01347_)
  );
  sg13g2_a22oi_1 _11697_ (
    .A1(_01325_),
    .A2(_01335_),
    .B1(_00109_),
    .B2(_01347_),
    .Y(_01348_)
  );
  sg13g2_nor4_1 _11698_ (
    .A(_00513_),
    .B(_01239_),
    .C(_01316_),
    .D(_01348_),
    .Y(_01349_)
  );
  sg13g2_buf_1 _11699_ (
    .A(_00215_),
    .X(_01350_)
  );
  sg13g2_nand3b_1 _11700_ (
    .A_N(addr_i_5_),
    .B(addr_i_6_),
    .C(addr_i_2_),
    .Y(_01352_)
  );
  sg13g2_buf_1 _11701_ (
    .A(_01352_),
    .X(_01353_)
  );
  sg13g2_buf_1 _11702_ (
    .A(_01353_),
    .X(_01354_)
  );
  sg13g2_buf_1 _11703_ (
    .A(_00828_),
    .X(_01355_)
  );
  sg13g2_a22oi_1 _11704_ (
    .A1(_01354_),
    .A2(_03391_),
    .B1(_01355_),
    .B2(_05834_),
    .Y(_01356_)
  );
  sg13g2_nor2_1 _11705_ (
    .A(addr_i_7_),
    .B(_01309_),
    .Y(_01357_)
  );
  sg13g2_or2_1 _11706_ (
    .A(_01356_),
    .B(_01357_),
    .X(_01358_)
  );
  sg13g2_nand2_1 _11707_ (
    .A(addr_i_12_),
    .B(addr_i_11_),
    .Y(_01359_)
  );
  sg13g2_nor2_1 _11708_ (
    .A(_07514_),
    .B(_01355_),
    .Y(_01360_)
  );
  sg13g2_nand3_1 _11709_ (
    .A(addr_i_5_),
    .B(_00802_),
    .C(_00290_),
    .Y(_01361_)
  );
  sg13g2_o21ai_1 _11710_ (
    .A1(addr_i_5_),
    .A2(_00440_),
    .B1(_01361_),
    .Y(_01363_)
  );
  sg13g2_nand2b_1 _11711_ (
    .A_N(_01360_),
    .B(_01363_),
    .Y(_01364_)
  );
  sg13g2_buf_1 _11712_ (
    .A(_00818_),
    .X(_01365_)
  );
  sg13g2_o21ai_1 _11713_ (
    .A1(_07547_),
    .A2(_01365_),
    .B1(addr_i_3_),
    .Y(_01366_)
  );
  sg13g2_buf_1 _11714_ (
    .A(_09393_),
    .X(_01367_)
  );
  sg13g2_nand2_1 _11715_ (
    .A(_05700_),
    .B(_04860_),
    .Y(_01368_)
  );
  sg13g2_nand2_1 _11716_ (
    .A(_01367_),
    .B(_01368_),
    .Y(_01369_)
  );
  sg13g2_nand3_1 _11717_ (
    .A(addr_i_4_),
    .B(_00581_),
    .C(_02020_),
    .Y(_01370_)
  );
  sg13g2_o21ai_1 _11718_ (
    .A1(addr_i_4_),
    .A2(_01369_),
    .B1(_01370_),
    .Y(_01371_)
  );
  sg13g2_a21oi_1 _11719_ (
    .A1(_01366_),
    .A2(_01371_),
    .B1(_03062_),
    .Y(_01372_)
  );
  sg13g2_nor2_1 _11720_ (
    .A(addr_i_9_),
    .B(_00201_),
    .Y(_01374_)
  );
  sg13g2_a21oi_1 _11721_ (
    .A1(addr_i_2_),
    .A2(addr_i_5_),
    .B1(addr_i_4_),
    .Y(_01375_)
  );
  sg13g2_nor2_1 _11722_ (
    .A(_00059_),
    .B(_01375_),
    .Y(_01376_)
  );
  sg13g2_nor3_1 _11723_ (
    .A(addr_i_5_),
    .B(_01019_),
    .C(_00542_),
    .Y(_01377_)
  );
  sg13g2_nor2_1 _11724_ (
    .A(addr_i_6_),
    .B(_07603_),
    .Y(_01378_)
  );
  sg13g2_o21ai_1 _11725_ (
    .A1(_01376_),
    .A2(_01377_),
    .B1(_01378_),
    .Y(_01379_)
  );
  sg13g2_buf_1 _11726_ (
    .A(_01106_),
    .X(_01380_)
  );
  sg13g2_a22oi_1 _11727_ (
    .A1(addr_i_3_),
    .A2(_00464_),
    .B1(_00346_),
    .B2(_01380_),
    .Y(_01381_)
  );
  sg13g2_nor2_1 _11728_ (
    .A(_06607_),
    .B(_07591_),
    .Y(_01382_)
  );
  sg13g2_nand2b_1 _11729_ (
    .A_N(_01381_),
    .B(_01382_),
    .Y(_01383_)
  );
  sg13g2_nand3_1 _11730_ (
    .A(_01374_),
    .B(_01379_),
    .C(_01383_),
    .Y(_01385_)
  );
  sg13g2_nand2_1 _11731_ (
    .A(addr_i_4_),
    .B(_08774_),
    .Y(_01386_)
  );
  sg13g2_nor2_1 _11732_ (
    .A(_01570_),
    .B(_06032_),
    .Y(_01387_)
  );
  sg13g2_nor2_1 _11733_ (
    .A(addr_i_3_),
    .B(_01387_),
    .Y(_01388_)
  );
  sg13g2_nand2_1 _11734_ (
    .A(addr_i_3_),
    .B(_01834_),
    .Y(_01389_)
  );
  sg13g2_nor2_1 _11735_ (
    .A(_03555_),
    .B(_01389_),
    .Y(_01390_)
  );
  sg13g2_buf_1 _11736_ (
    .A(_08674_),
    .X(_01391_)
  );
  sg13g2_a22oi_1 _11737_ (
    .A1(_01386_),
    .A2(_01388_),
    .B1(_01390_),
    .B2(_01391_),
    .Y(_01392_)
  );
  sg13g2_nor3_1 _11738_ (
    .A(_01372_),
    .B(_01385_),
    .C(_01392_),
    .Y(_01393_)
  );
  sg13g2_a22oi_1 _11739_ (
    .A1(addr_i_9_),
    .A2(_01364_),
    .B1(_01393_),
    .B2(addr_i_10_),
    .Y(_01394_)
  );
  sg13g2_a22oi_1 _11740_ (
    .A1(_01350_),
    .A2(_01358_),
    .B1(_01359_),
    .B2(_01394_),
    .Y(_01396_)
  );
  sg13g2_o21ai_1 _11741_ (
    .A1(_03621_),
    .A2(_03523_),
    .B1(_08156_),
    .Y(_01397_)
  );
  sg13g2_nand2_1 _11742_ (
    .A(addr_i_3_),
    .B(_07237_),
    .Y(_01398_)
  );
  sg13g2_and2_1 _11743_ (
    .A(_01397_),
    .B(_01398_),
    .X(_01399_)
  );
  sg13g2_nor2_1 _11744_ (
    .A(_06375_),
    .B(_00972_),
    .Y(_01400_)
  );
  sg13g2_nor2_1 _11745_ (
    .A(_07933_),
    .B(_00198_),
    .Y(_01401_)
  );
  sg13g2_buf_1 _11746_ (
    .A(_01401_),
    .X(_01402_)
  );
  sg13g2_a22oi_1 _11747_ (
    .A1(addr_i_3_),
    .A2(_01400_),
    .B1(_01402_),
    .B2(addr_i_2_),
    .Y(_01403_)
  );
  sg13g2_a22oi_1 _11748_ (
    .A1(addr_i_2_),
    .A2(_01399_),
    .B1(_01403_),
    .B2(_08487_),
    .Y(_01404_)
  );
  sg13g2_nor3_1 _11749_ (
    .A(_08045_),
    .B(_02613_),
    .C(_02843_),
    .Y(_01405_)
  );
  sg13g2_nor3_1 _11750_ (
    .A(addr_i_7_),
    .B(addr_i_5_),
    .C(_07812_),
    .Y(_01407_)
  );
  sg13g2_nor2_1 _11751_ (
    .A(_02196_),
    .B(_01228_),
    .Y(_01408_)
  );
  sg13g2_o21ai_1 _11752_ (
    .A1(_01407_),
    .A2(_01408_),
    .B1(addr_i_6_),
    .Y(_01409_)
  );
  sg13g2_nand2_1 _11753_ (
    .A(_07061_),
    .B(_03172_),
    .Y(_01410_)
  );
  sg13g2_o21ai_1 _11754_ (
    .A1(_00597_),
    .A2(_00632_),
    .B1(addr_i_3_),
    .Y(_01411_)
  );
  sg13g2_nand3_1 _11755_ (
    .A(_01409_),
    .B(_01410_),
    .C(_01411_),
    .Y(_01412_)
  );
  sg13g2_nor2_1 _11756_ (
    .A(addr_i_7_),
    .B(_06099_),
    .Y(_01413_)
  );
  sg13g2_nand2_1 _11757_ (
    .A(_08100_),
    .B(_00442_),
    .Y(_01414_)
  );
  sg13g2_a21oi_1 _11758_ (
    .A1(_04229_),
    .A2(_01414_),
    .B1(addr_i_6_),
    .Y(_01415_)
  );
  sg13g2_a221oi_1 _11759_ (
    .A1(addr_i_4_),
    .A2(_01412_),
    .B1(_01413_),
    .B2(_01202_),
    .C1(_01415_),
    .Y(_01416_)
  );
  sg13g2_nor2_1 _11760_ (
    .A(addr_i_8_),
    .B(_01416_),
    .Y(_01418_)
  );
  sg13g2_nor3_1 _11761_ (
    .A(_01404_),
    .B(_01405_),
    .C(_01418_),
    .Y(_01419_)
  );
  sg13g2_buf_1 _11762_ (
    .A(_03194_),
    .X(_01420_)
  );
  sg13g2_nor2_1 _11763_ (
    .A(addr_i_7_),
    .B(_00557_),
    .Y(_01421_)
  );
  sg13g2_nand2_1 _11764_ (
    .A(_04362_),
    .B(_01976_),
    .Y(_01422_)
  );
  sg13g2_a221oi_1 _11765_ (
    .A1(_01420_),
    .A2(_01421_),
    .B1(_01422_),
    .B2(_01262_),
    .C1(_00116_),
    .Y(_01423_)
  );
  sg13g2_nor2_1 _11766_ (
    .A(_01373_),
    .B(_02558_),
    .Y(_01424_)
  );
  sg13g2_nand2_1 _11767_ (
    .A(_05390_),
    .B(_05424_),
    .Y(_01425_)
  );
  sg13g2_a21oi_1 _11768_ (
    .A1(_00907_),
    .A2(_01425_),
    .B1(_06619_),
    .Y(_01426_)
  );
  sg13g2_nor3_1 _11769_ (
    .A(_00105_),
    .B(_00159_),
    .C(_04915_),
    .Y(_01427_)
  );
  sg13g2_nor4_1 _11770_ (
    .A(addr_i_3_),
    .B(_01424_),
    .C(_01426_),
    .D(_01427_),
    .Y(_01429_)
  );
  sg13g2_a21oi_1 _11771_ (
    .A1(_09474_),
    .A2(_01216_),
    .B1(addr_i_8_),
    .Y(_01430_)
  );
  sg13g2_o21ai_1 _11772_ (
    .A1(_01423_),
    .A2(_01429_),
    .B1(_01430_),
    .Y(_01431_)
  );
  sg13g2_buf_1 _11773_ (
    .A(_01406_),
    .X(_01432_)
  );
  sg13g2_nand2_1 _11774_ (
    .A(_04285_),
    .B(_01432_),
    .Y(_01433_)
  );
  sg13g2_a21oi_1 _11775_ (
    .A1(_02349_),
    .A2(_00404_),
    .B1(addr_i_4_),
    .Y(_01434_)
  );
  sg13g2_a22oi_1 _11776_ (
    .A1(addr_i_4_),
    .A2(_01433_),
    .B1(_01434_),
    .B2(_00026_),
    .Y(_01435_)
  );
  sg13g2_buf_1 _11777_ (
    .A(_03106_),
    .X(_01436_)
  );
  sg13g2_nand2_1 _11778_ (
    .A(_08376_),
    .B(_00678_),
    .Y(_01437_)
  );
  sg13g2_or3_1 _11779_ (
    .A(addr_i_4_),
    .B(addr_i_7_),
    .C(addr_i_6_),
    .X(_01438_)
  );
  sg13g2_o21ai_1 _11780_ (
    .A1(_01436_),
    .A2(_01437_),
    .B1(_01438_),
    .Y(_01440_)
  );
  sg13g2_buf_1 _11781_ (
    .A(_00680_),
    .X(_01441_)
  );
  sg13g2_a21oi_1 _11782_ (
    .A1(_01065_),
    .A2(_01441_),
    .B1(_01252_),
    .Y(_01442_)
  );
  sg13g2_a22oi_1 _11783_ (
    .A1(addr_i_2_),
    .A2(_01440_),
    .B1(_01442_),
    .B2(_04506_),
    .Y(_01443_)
  );
  sg13g2_mux2_1 _11784_ (
    .A0(_01435_),
    .A1(_01443_),
    .S(_01169_),
    .X(_01444_)
  );
  sg13g2_buf_1 _11785_ (
    .A(_04528_),
    .X(_01445_)
  );
  sg13g2_nand2_1 _11786_ (
    .A(_01445_),
    .B(_00209_),
    .Y(_01446_)
  );
  sg13g2_nand3_1 _11787_ (
    .A(addr_i_8_),
    .B(_01444_),
    .C(_01446_),
    .Y(_01447_)
  );
  sg13g2_nand3_1 _11788_ (
    .A(_01176_),
    .B(_01431_),
    .C(_01447_),
    .Y(_01448_)
  );
  sg13g2_o21ai_1 _11789_ (
    .A1(_00109_),
    .A2(_01419_),
    .B1(_01448_),
    .Y(_01449_)
  );
  sg13g2_nand2_1 _11790_ (
    .A(addr_i_12_),
    .B(_03029_),
    .Y(_01451_)
  );
  sg13g2_nand2_1 _11791_ (
    .A(_03731_),
    .B(addr_i_9_),
    .Y(_01452_)
  );
  sg13g2_nand2_1 _11792_ (
    .A(_00593_),
    .B(_09493_),
    .Y(_01453_)
  );
  sg13g2_a21oi_1 _11793_ (
    .A1(_01453_),
    .A2(_01398_),
    .B1(_01343_),
    .Y(_01454_)
  );
  sg13g2_o21ai_1 _11794_ (
    .A1(_07911_),
    .A2(_00660_),
    .B1(addr_i_8_),
    .Y(_01455_)
  );
  sg13g2_nor2_1 _11795_ (
    .A(_00020_),
    .B(_02733_),
    .Y(_01456_)
  );
  sg13g2_a21oi_1 _11796_ (
    .A1(_01336_),
    .A2(_00844_),
    .B1(_01456_),
    .Y(_01457_)
  );
  sg13g2_nor2_1 _11797_ (
    .A(_00390_),
    .B(_01457_),
    .Y(_01458_)
  );
  sg13g2_buf_1 _11798_ (
    .A(_08885_),
    .X(_01459_)
  );
  sg13g2_nand2_1 _11799_ (
    .A(_01459_),
    .B(_00960_),
    .Y(_01460_)
  );
  sg13g2_nand2_1 _11800_ (
    .A(addr_i_3_),
    .B(_03194_),
    .Y(_01462_)
  );
  sg13g2_nand2_1 _11801_ (
    .A(_05845_),
    .B(_00768_),
    .Y(_01463_)
  );
  sg13g2_nand2_1 _11802_ (
    .A(_01462_),
    .B(_01463_),
    .Y(_01464_)
  );
  sg13g2_nand2_1 _11803_ (
    .A(addr_i_5_),
    .B(_01464_),
    .Y(_01465_)
  );
  sg13g2_a21oi_1 _11804_ (
    .A1(_01460_),
    .A2(_01465_),
    .B1(_00507_),
    .Y(_01466_)
  );
  sg13g2_nor4_1 _11805_ (
    .A(_01454_),
    .B(_01455_),
    .C(_01458_),
    .D(_01466_),
    .Y(_01467_)
  );
  sg13g2_o21ai_1 _11806_ (
    .A1(_01070_),
    .A2(_02744_),
    .B1(_00250_),
    .Y(_01468_)
  );
  sg13g2_a21oi_1 _11807_ (
    .A1(_00070_),
    .A2(_00105_),
    .B1(_01339_),
    .Y(_01469_)
  );
  sg13g2_a21oi_1 _11808_ (
    .A1(_03292_),
    .A2(_01468_),
    .B1(_01469_),
    .Y(_01470_)
  );
  sg13g2_nor2_1 _11809_ (
    .A(addr_i_3_),
    .B(_06873_),
    .Y(_01471_)
  );
  sg13g2_buf_1 _11810_ (
    .A(_02602_),
    .X(_01473_)
  );
  sg13g2_a21oi_1 _11811_ (
    .A1(_01473_),
    .A2(_00339_),
    .B1(_00726_),
    .Y(_01474_)
  );
  sg13g2_buf_1 _11812_ (
    .A(_03820_),
    .X(_01475_)
  );
  sg13g2_o21ai_1 _11813_ (
    .A1(_01471_),
    .A2(_01474_),
    .B1(_01475_),
    .Y(_01476_)
  );
  sg13g2_a21oi_1 _11814_ (
    .A1(_01470_),
    .A2(_01476_),
    .B1(addr_i_6_),
    .Y(_01477_)
  );
  sg13g2_nor2_1 _11815_ (
    .A(_05856_),
    .B(_01179_),
    .Y(_01478_)
  );
  sg13g2_nor3_1 _11816_ (
    .A(_00053_),
    .B(_01375_),
    .C(_01478_),
    .Y(_01479_)
  );
  sg13g2_buf_1 _11817_ (
    .A(_01244_),
    .X(_01480_)
  );
  sg13g2_buf_1 _11818_ (
    .A(_02294_),
    .X(_01481_)
  );
  sg13g2_a22oi_1 _11819_ (
    .A1(_00467_),
    .A2(_02536_),
    .B1(_01480_),
    .B2(_01481_),
    .Y(_01482_)
  );
  sg13g2_nor4_1 _11820_ (
    .A(addr_i_8_),
    .B(_01477_),
    .C(_01479_),
    .D(_01482_),
    .Y(_01484_)
  );
  sg13g2_nor3_1 _11821_ (
    .A(_01452_),
    .B(_01467_),
    .C(_01484_),
    .Y(_01485_)
  );
  sg13g2_nor2_1 _11822_ (
    .A(addr_i_6_),
    .B(_04926_),
    .Y(_01486_)
  );
  sg13g2_nor2_1 _11823_ (
    .A(addr_i_4_),
    .B(_01486_),
    .Y(_01487_)
  );
  sg13g2_a21oi_1 _11824_ (
    .A1(_09474_),
    .A2(_01365_),
    .B1(_01487_),
    .Y(_01488_)
  );
  sg13g2_nor3_1 _11825_ (
    .A(_03930_),
    .B(addr_i_6_),
    .C(_05833_),
    .Y(_01489_)
  );
  sg13g2_o21ai_1 _11826_ (
    .A1(_00023_),
    .A2(_01489_),
    .B1(addr_i_4_),
    .Y(_01490_)
  );
  sg13g2_o21ai_1 _11827_ (
    .A1(addr_i_5_),
    .A2(_01488_),
    .B1(_01490_),
    .Y(_01491_)
  );
  sg13g2_nand2_1 _11828_ (
    .A(addr_i_3_),
    .B(_01491_),
    .Y(_01492_)
  );
  sg13g2_nand2_1 _11829_ (
    .A(_04418_),
    .B(_00863_),
    .Y(_01493_)
  );
  sg13g2_nor2_1 _11830_ (
    .A(_08100_),
    .B(_00086_),
    .Y(_01495_)
  );
  sg13g2_o21ai_1 _11831_ (
    .A1(_07625_),
    .A2(_01495_),
    .B1(_01691_),
    .Y(_01496_)
  );
  sg13g2_nand2_1 _11832_ (
    .A(addr_i_8_),
    .B(_00131_),
    .Y(_01497_)
  );
  sg13g2_a221oi_1 _11833_ (
    .A1(addr_i_7_),
    .A2(_01493_),
    .B1(_01496_),
    .B2(_00048_),
    .C1(_01497_),
    .Y(_01498_)
  );
  sg13g2_buf_1 _11834_ (
    .A(_01222_),
    .X(_01499_)
  );
  sg13g2_buf_1 _11835_ (
    .A(_01014_),
    .X(_01500_)
  );
  sg13g2_o21ai_1 _11836_ (
    .A1(_01262_),
    .A2(_01500_),
    .B1(addr_i_3_),
    .Y(_01501_)
  );
  sg13g2_nand3_1 _11837_ (
    .A(_05357_),
    .B(_01499_),
    .C(_01501_),
    .Y(_01502_)
  );
  sg13g2_o21ai_1 _11838_ (
    .A1(_07712_),
    .A2(_00436_),
    .B1(addr_i_3_),
    .Y(_01503_)
  );
  sg13g2_nand2_1 _11839_ (
    .A(_01319_),
    .B(_00819_),
    .Y(_01504_)
  );
  sg13g2_nand3_1 _11840_ (
    .A(_06706_),
    .B(_01503_),
    .C(_01504_),
    .Y(_01506_)
  );
  sg13g2_buf_1 _11841_ (
    .A(_04926_),
    .X(_01507_)
  );
  sg13g2_buf_1 _11842_ (
    .A(_01507_),
    .X(_01508_)
  );
  sg13g2_nor3_1 _11843_ (
    .A(addr_i_3_),
    .B(_01508_),
    .C(_01380_),
    .Y(_01509_)
  );
  sg13g2_a22oi_1 _11844_ (
    .A1(addr_i_3_),
    .A2(_00747_),
    .B1(_01509_),
    .B2(addr_i_6_),
    .Y(_01510_)
  );
  sg13g2_a22oi_1 _11845_ (
    .A1(addr_i_4_),
    .A2(_01502_),
    .B1(_01506_),
    .B2(_01510_),
    .Y(_01511_)
  );
  sg13g2_a22oi_1 _11846_ (
    .A1(_01492_),
    .A2(_01498_),
    .B1(_01511_),
    .B2(_00774_),
    .Y(_01512_)
  );
  sg13g2_nor4_1 _11847_ (
    .A(_01449_),
    .B(_01451_),
    .C(_01485_),
    .D(_01512_),
    .Y(_01513_)
  );
  sg13g2_nor4_1 _11848_ (
    .A(_01210_),
    .B(_01349_),
    .C(_01396_),
    .D(_01513_),
    .Y(data_o_12_)
  );
  sg13g2_buf_1 _11849_ (
    .A(_03732_),
    .X(_01514_)
  );
  sg13g2_o21ai_1 _11850_ (
    .A1(_07889_),
    .A2(_01514_),
    .B1(_02898_),
    .Y(_01516_)
  );
  sg13g2_buf_1 _11851_ (
    .A(_08332_),
    .X(_01517_)
  );
  sg13g2_nor2_1 _11852_ (
    .A(_01517_),
    .B(_00213_),
    .Y(_01518_)
  );
  sg13g2_buf_1 _11853_ (
    .A(_05379_),
    .X(_01519_)
  );
  sg13g2_buf_1 _11854_ (
    .A(_04373_),
    .X(_01520_)
  );
  sg13g2_o21ai_1 _11855_ (
    .A1(_01282_),
    .A2(_01519_),
    .B1(_01520_),
    .Y(_01521_)
  );
  sg13g2_nand3_1 _11856_ (
    .A(_00353_),
    .B(_01518_),
    .C(_01521_),
    .Y(_01522_)
  );
  sg13g2_a221oi_1 _11857_ (
    .A1(_00626_),
    .A2(_01305_),
    .B1(_01516_),
    .B2(addr_i_2_),
    .C1(_01522_),
    .Y(_01523_)
  );
  sg13g2_nand2_1 _11858_ (
    .A(_09038_),
    .B(_00664_),
    .Y(_01524_)
  );
  sg13g2_a21o_1 _11859_ (
    .A1(_00943_),
    .A2(_01524_),
    .B1(_08000_),
    .X(_01525_)
  );
  sg13g2_buf_1 _11860_ (
    .A(_00725_),
    .X(_01527_)
  );
  sg13g2_buf_1 _11861_ (
    .A(_01113_),
    .X(_01528_)
  );
  sg13g2_a21oi_1 _11862_ (
    .A1(_01527_),
    .A2(_01450_),
    .B1(_01528_),
    .Y(_01529_)
  );
  sg13g2_nor2_1 _11863_ (
    .A(addr_i_2_),
    .B(_08609_),
    .Y(_01530_)
  );
  sg13g2_a22oi_1 _11864_ (
    .A1(addr_i_3_),
    .A2(_04727_),
    .B1(_01530_),
    .B2(addr_i_4_),
    .Y(_01531_)
  );
  sg13g2_a21oi_1 _11865_ (
    .A1(_01525_),
    .A2(_01529_),
    .B1(_01531_),
    .Y(_01532_)
  );
  sg13g2_o21ai_1 _11866_ (
    .A1(_06264_),
    .A2(_01049_),
    .B1(addr_i_3_),
    .Y(_01533_)
  );
  sg13g2_a21oi_1 _11867_ (
    .A1(_03391_),
    .A2(_01533_),
    .B1(addr_i_7_),
    .Y(_01534_)
  );
  sg13g2_a22oi_1 _11868_ (
    .A1(addr_i_7_),
    .A2(_01532_),
    .B1(_01534_),
    .B2(addr_i_8_),
    .Y(_01535_)
  );
  sg13g2_a21oi_1 _11869_ (
    .A1(_01462_),
    .A2(_01463_),
    .B1(addr_i_5_),
    .Y(_01536_)
  );
  sg13g2_a21oi_1 _11870_ (
    .A1(_00703_),
    .A2(_00401_),
    .B1(_01536_),
    .Y(_01538_)
  );
  sg13g2_a21oi_1 _11871_ (
    .A1(addr_i_4_),
    .A2(addr_i_5_),
    .B1(addr_i_2_),
    .Y(_01539_)
  );
  sg13g2_a21oi_1 _11872_ (
    .A1(_00650_),
    .A2(_05689_),
    .B1(addr_i_3_),
    .Y(_01540_)
  );
  sg13g2_a21o_1 _11873_ (
    .A1(addr_i_3_),
    .A2(_01539_),
    .B1(_01540_),
    .X(_01541_)
  );
  sg13g2_buf_1 _11874_ (
    .A(_01867_),
    .X(_01542_)
  );
  sg13g2_buf_1 _11875_ (
    .A(_02371_),
    .X(_01543_)
  );
  sg13g2_nand2_1 _11876_ (
    .A(_00158_),
    .B(_08111_),
    .Y(_01544_)
  );
  sg13g2_o21ai_1 _11877_ (
    .A1(_01543_),
    .A2(_01544_),
    .B1(addr_i_8_),
    .Y(_01545_)
  );
  sg13g2_a221oi_1 _11878_ (
    .A1(_00466_),
    .A2(_00872_),
    .B1(_01541_),
    .B2(_01542_),
    .C1(_01545_),
    .Y(_01546_)
  );
  sg13g2_o21ai_1 _11879_ (
    .A1(_00507_),
    .A2(_01538_),
    .B1(_01546_),
    .Y(_01547_)
  );
  sg13g2_nand3b_1 _11880_ (
    .A_N(_01535_),
    .B(_01547_),
    .C(addr_i_9_),
    .Y(_01549_)
  );
  sg13g2_nand3b_1 _11881_ (
    .A_N(_01523_),
    .B(addr_i_10_),
    .C(_01549_),
    .Y(_01550_)
  );
  sg13g2_nor2_1 _11882_ (
    .A(addr_i_3_),
    .B(_01603_),
    .Y(_01551_)
  );
  sg13g2_nor2_1 _11883_ (
    .A(_01965_),
    .B(_08941_),
    .Y(_01552_)
  );
  sg13g2_o21ai_1 _11884_ (
    .A1(_01551_),
    .A2(_01552_),
    .B1(_06154_),
    .Y(_01553_)
  );
  sg13g2_nand2_1 _11885_ (
    .A(_00006_),
    .B(_00736_),
    .Y(_01554_)
  );
  sg13g2_nand2_1 _11886_ (
    .A(addr_i_6_),
    .B(_02459_),
    .Y(_01555_)
  );
  sg13g2_a21oi_1 _11887_ (
    .A1(_00650_),
    .A2(_01555_),
    .B1(_05070_),
    .Y(_01556_)
  );
  sg13g2_a22oi_1 _11888_ (
    .A1(_04373_),
    .A2(_01554_),
    .B1(_01556_),
    .B2(addr_i_8_),
    .Y(_01557_)
  );
  sg13g2_nand2_1 _11889_ (
    .A(_01553_),
    .B(_01557_),
    .Y(_01558_)
  );
  sg13g2_nor2_1 _11890_ (
    .A(addr_i_4_),
    .B(_00016_),
    .Y(_01560_)
  );
  sg13g2_o21ai_1 _11891_ (
    .A1(_00226_),
    .A2(_01560_),
    .B1(addr_i_3_),
    .Y(_01561_)
  );
  sg13g2_o21ai_1 _11892_ (
    .A1(_07812_),
    .A2(_00110_),
    .B1(addr_i_5_),
    .Y(_01562_)
  );
  sg13g2_a21oi_1 _11893_ (
    .A1(_01561_),
    .A2(_01562_),
    .B1(addr_i_6_),
    .Y(_01563_)
  );
  sg13g2_o21ai_1 _11894_ (
    .A1(_01558_),
    .A2(_01563_),
    .B1(_09315_),
    .Y(_01564_)
  );
  sg13g2_a21oi_1 _11895_ (
    .A1(_09492_),
    .A2(_01439_),
    .B1(_00792_),
    .Y(_01565_)
  );
  sg13g2_o21ai_1 _11896_ (
    .A1(addr_i_5_),
    .A2(_01565_),
    .B1(_06784_),
    .Y(_01566_)
  );
  sg13g2_nor2_1 _11897_ (
    .A(addr_i_4_),
    .B(_04561_),
    .Y(_01567_)
  );
  sg13g2_a21oi_1 _11898_ (
    .A1(_02218_),
    .A2(_01368_),
    .B1(_09492_),
    .Y(_01568_)
  );
  sg13g2_nor2_1 _11899_ (
    .A(_01567_),
    .B(_01568_),
    .Y(_01569_)
  );
  sg13g2_buf_1 _11900_ (
    .A(_01244_),
    .X(_01571_)
  );
  sg13g2_nand2_1 _11901_ (
    .A(addr_i_6_),
    .B(_00964_),
    .Y(_01572_)
  );
  sg13g2_a22oi_1 _11902_ (
    .A1(_01571_),
    .A2(_01572_),
    .B1(addr_i_2_),
    .B2(_09502_),
    .Y(_01573_)
  );
  sg13g2_a21oi_1 _11903_ (
    .A1(addr_i_2_),
    .A2(_01569_),
    .B1(_01573_),
    .Y(_01574_)
  );
  sg13g2_o21ai_1 _11904_ (
    .A1(_01566_),
    .A2(_01574_),
    .B1(addr_i_8_),
    .Y(_01575_)
  );
  sg13g2_nand2b_1 _11905_ (
    .A_N(_01564_),
    .B(_01575_),
    .Y(_01576_)
  );
  sg13g2_nor2_1 _11906_ (
    .A(_00246_),
    .B(_00521_),
    .Y(_01577_)
  );
  sg13g2_a22oi_1 _11907_ (
    .A1(addr_i_3_),
    .A2(_00110_),
    .B1(_00667_),
    .B2(_01577_),
    .Y(_01578_)
  );
  sg13g2_nor2_1 _11908_ (
    .A(_07049_),
    .B(_03798_),
    .Y(_01579_)
  );
  sg13g2_buf_1 _11909_ (
    .A(_01579_),
    .X(_01580_)
  );
  sg13g2_nor2_1 _11910_ (
    .A(_05734_),
    .B(_07469_),
    .Y(_01582_)
  );
  sg13g2_a21oi_1 _11911_ (
    .A1(_01580_),
    .A2(_01275_),
    .B1(_01582_),
    .Y(_01583_)
  );
  sg13g2_o21ai_1 _11912_ (
    .A1(addr_i_6_),
    .A2(_01578_),
    .B1(_01583_),
    .Y(_01584_)
  );
  sg13g2_buf_1 _11913_ (
    .A(_09050_),
    .X(_01585_)
  );
  sg13g2_nand2_1 _11914_ (
    .A(_01585_),
    .B(_00244_),
    .Y(_01586_)
  );
  sg13g2_buf_1 _11915_ (
    .A(_00154_),
    .X(_01587_)
  );
  sg13g2_buf_1 _11916_ (
    .A(_03303_),
    .X(_01588_)
  );
  sg13g2_nand3_1 _11917_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .C(addr_i_6_),
    .Y(_01589_)
  );
  sg13g2_nand2_1 _11918_ (
    .A(_01588_),
    .B(_01589_),
    .Y(_01590_)
  );
  sg13g2_nand2_1 _11919_ (
    .A(_01587_),
    .B(_01590_),
    .Y(_01591_)
  );
  sg13g2_a21oi_1 _11920_ (
    .A1(_01586_),
    .A2(_01591_),
    .B1(addr_i_3_),
    .Y(_01593_)
  );
  sg13g2_nand2_1 _11921_ (
    .A(_00292_),
    .B(_07248_),
    .Y(_01594_)
  );
  sg13g2_nand2_1 _11922_ (
    .A(addr_i_8_),
    .B(_01594_),
    .Y(_01595_)
  );
  sg13g2_a22oi_1 _11923_ (
    .A1(_01279_),
    .A2(_01584_),
    .B1(_01593_),
    .B2(_01595_),
    .Y(_01596_)
  );
  sg13g2_a21oi_1 _11924_ (
    .A1(addr_i_7_),
    .A2(_02218_),
    .B1(_09393_),
    .Y(_01597_)
  );
  sg13g2_a21oi_1 _11925_ (
    .A1(_00547_),
    .A2(_00763_),
    .B1(addr_i_3_),
    .Y(_01598_)
  );
  sg13g2_a22oi_1 _11926_ (
    .A1(_00783_),
    .A2(_01294_),
    .B1(_01597_),
    .B2(_01598_),
    .Y(_01599_)
  );
  sg13g2_inv_1 _11927_ (
    .A(_01599_),
    .Y(_01600_)
  );
  sg13g2_nand2_1 _11928_ (
    .A(_08089_),
    .B(_04860_),
    .Y(_01601_)
  );
  sg13g2_and2_1 _11929_ (
    .A(_00763_),
    .B(_01601_),
    .X(_01602_)
  );
  sg13g2_nor2_1 _11930_ (
    .A(_00246_),
    .B(_02020_),
    .Y(_01604_)
  );
  sg13g2_a22oi_1 _11931_ (
    .A1(addr_i_2_),
    .A2(_01228_),
    .B1(_01604_),
    .B2(_09508_),
    .Y(_01605_)
  );
  sg13g2_a22oi_1 _11932_ (
    .A1(addr_i_3_),
    .A2(_01602_),
    .B1(_01605_),
    .B2(addr_i_4_),
    .Y(_01606_)
  );
  sg13g2_a22oi_1 _11933_ (
    .A1(addr_i_4_),
    .A2(_01600_),
    .B1(_01606_),
    .B2(addr_i_8_),
    .Y(_01607_)
  );
  sg13g2_o21ai_1 _11934_ (
    .A1(_01596_),
    .A2(_01607_),
    .B1(addr_i_9_),
    .Y(_01608_)
  );
  sg13g2_a21o_1 _11935_ (
    .A1(_01576_),
    .A2(_01608_),
    .B1(addr_i_10_),
    .X(_01609_)
  );
  sg13g2_nand2_1 _11936_ (
    .A(_00374_),
    .B(addr_i_8_),
    .Y(_01610_)
  );
  sg13g2_buf_1 _11937_ (
    .A(_01610_),
    .X(_01611_)
  );
  sg13g2_buf_1 _11938_ (
    .A(_01611_),
    .X(_01612_)
  );
  sg13g2_nor2_1 _11939_ (
    .A(_03731_),
    .B(_01612_),
    .Y(_01613_)
  );
  sg13g2_buf_1 _11940_ (
    .A(_08332_),
    .X(_01615_)
  );
  sg13g2_buf_1 _11941_ (
    .A(_00557_),
    .X(_01616_)
  );
  sg13g2_o21ai_1 _11942_ (
    .A1(_01615_),
    .A2(_01616_),
    .B1(_08011_),
    .Y(_01617_)
  );
  sg13g2_nand2_1 _11943_ (
    .A(_00294_),
    .B(_00011_),
    .Y(_01618_)
  );
  sg13g2_nand3_1 _11944_ (
    .A(_00390_),
    .B(_01617_),
    .C(_01618_),
    .Y(_01619_)
  );
  sg13g2_a21oi_1 _11945_ (
    .A1(_01354_),
    .A2(_01199_),
    .B1(addr_i_4_),
    .Y(_01620_)
  );
  sg13g2_a22oi_1 _11946_ (
    .A1(addr_i_4_),
    .A2(_01619_),
    .B1(_01620_),
    .B2(_00048_),
    .Y(_01621_)
  );
  sg13g2_nand2_1 _11947_ (
    .A(addr_i_7_),
    .B(_06077_),
    .Y(_01622_)
  );
  sg13g2_nor2_1 _11948_ (
    .A(addr_i_2_),
    .B(_01622_),
    .Y(_01623_)
  );
  sg13g2_o21ai_1 _11949_ (
    .A1(addr_i_7_),
    .A2(_08553_),
    .B1(_00371_),
    .Y(_01624_)
  );
  sg13g2_a221oi_1 _11950_ (
    .A1(addr_i_4_),
    .A2(_01623_),
    .B1(_01624_),
    .B2(addr_i_2_),
    .C1(addr_i_3_),
    .Y(_01626_)
  );
  sg13g2_nor2_1 _11951_ (
    .A(_00019_),
    .B(_07160_),
    .Y(_01627_)
  );
  sg13g2_nor2_1 _11952_ (
    .A(_00550_),
    .B(_01276_),
    .Y(_01628_)
  );
  sg13g2_nor2_1 _11953_ (
    .A(addr_i_7_),
    .B(_01628_),
    .Y(_01629_)
  );
  sg13g2_buf_1 _11954_ (
    .A(_00360_),
    .X(_01630_)
  );
  sg13g2_o21ai_1 _11955_ (
    .A1(_01627_),
    .A2(_01629_),
    .B1(_01630_),
    .Y(_01631_)
  );
  sg13g2_o21ai_1 _11956_ (
    .A1(_01621_),
    .A2(_01626_),
    .B1(_01631_),
    .Y(_01632_)
  );
  sg13g2_buf_1 _11957_ (
    .A(_00429_),
    .X(_01633_)
  );
  sg13g2_nand2_1 _11958_ (
    .A(_01174_),
    .B(_01633_),
    .Y(_01634_)
  );
  sg13g2_nor2_1 _11959_ (
    .A(_03128_),
    .B(_03512_),
    .Y(_01635_)
  );
  sg13g2_nor2_1 _11960_ (
    .A(addr_i_3_),
    .B(_03117_),
    .Y(_01637_)
  );
  sg13g2_a22oi_1 _11961_ (
    .A1(addr_i_3_),
    .A2(_01635_),
    .B1(_01637_),
    .B2(addr_i_2_),
    .Y(_01638_)
  );
  sg13g2_nor2_1 _11962_ (
    .A(_00518_),
    .B(_01638_),
    .Y(_01639_)
  );
  sg13g2_buf_1 _11963_ (
    .A(_03029_),
    .X(_01640_)
  );
  sg13g2_o21ai_1 _11964_ (
    .A1(_01634_),
    .A2(_01639_),
    .B1(_01640_),
    .Y(_01641_)
  );
  sg13g2_a221oi_1 _11965_ (
    .A1(_01550_),
    .A2(_01609_),
    .B1(_01613_),
    .B2(_01632_),
    .C1(_01641_),
    .Y(_01642_)
  );
  sg13g2_nor2_1 _11966_ (
    .A(_00034_),
    .B(_01353_),
    .Y(_01643_)
  );
  sg13g2_nand2_1 _11967_ (
    .A(addr_i_7_),
    .B(_03391_),
    .Y(_01644_)
  );
  sg13g2_nor2_1 _11968_ (
    .A(addr_i_7_),
    .B(_00008_),
    .Y(_01645_)
  );
  sg13g2_nor2_1 _11969_ (
    .A(_00807_),
    .B(_01645_),
    .Y(_01646_)
  );
  sg13g2_o21ai_1 _11970_ (
    .A1(_01643_),
    .A2(_01644_),
    .B1(_01646_),
    .Y(_01648_)
  );
  sg13g2_nand2_1 _11971_ (
    .A(addr_i_6_),
    .B(_08254_),
    .Y(_01649_)
  );
  sg13g2_a21oi_1 _11972_ (
    .A1(_01103_),
    .A2(_00762_),
    .B1(addr_i_4_),
    .Y(_01650_)
  );
  sg13g2_a22oi_1 _11973_ (
    .A1(addr_i_4_),
    .A2(_01649_),
    .B1(_01650_),
    .B2(_08674_),
    .Y(_01651_)
  );
  sg13g2_buf_1 _11974_ (
    .A(_00738_),
    .X(_01652_)
  );
  sg13g2_buf_1 _11975_ (
    .A(_01652_),
    .X(_01653_)
  );
  sg13g2_a21oi_1 _11976_ (
    .A1(addr_i_6_),
    .A2(_00380_),
    .B1(_05700_),
    .Y(_01654_)
  );
  sg13g2_o21ai_1 _11977_ (
    .A1(_01653_),
    .A2(_01654_),
    .B1(addr_i_2_),
    .Y(_01655_)
  );
  sg13g2_buf_1 _11978_ (
    .A(_00448_),
    .X(_01656_)
  );
  sg13g2_o21ai_1 _11979_ (
    .A1(_03227_),
    .A2(_01656_),
    .B1(_00385_),
    .Y(_01657_)
  );
  sg13g2_nor2_1 _11980_ (
    .A(_07933_),
    .B(_04064_),
    .Y(_01659_)
  );
  sg13g2_buf_1 _11981_ (
    .A(_01659_),
    .X(_01660_)
  );
  sg13g2_o21ai_1 _11982_ (
    .A1(_01660_),
    .A2(_01107_),
    .B1(addr_i_3_),
    .Y(_01661_)
  );
  sg13g2_a21o_1 _11983_ (
    .A1(_09483_),
    .A2(_09475_),
    .B1(addr_i_3_),
    .X(_01662_)
  );
  sg13g2_nand2_1 _11984_ (
    .A(addr_i_6_),
    .B(_00418_),
    .Y(_01663_)
  );
  sg13g2_a21oi_1 _11985_ (
    .A1(_01661_),
    .A2(_01662_),
    .B1(_01663_),
    .Y(_01664_)
  );
  sg13g2_a22oi_1 _11986_ (
    .A1(_01651_),
    .A2(_01655_),
    .B1(_01657_),
    .B2(_01664_),
    .Y(_01665_)
  );
  sg13g2_buf_1 _11987_ (
    .A(_01310_),
    .X(_01666_)
  );
  sg13g2_nand2_1 _11988_ (
    .A(_01666_),
    .B(_00844_),
    .Y(_01667_)
  );
  sg13g2_nand2_1 _11989_ (
    .A(_00588_),
    .B(_01656_),
    .Y(_01668_)
  );
  sg13g2_a21oi_1 _11990_ (
    .A1(_01667_),
    .A2(_01668_),
    .B1(_04705_),
    .Y(_01670_)
  );
  sg13g2_a22oi_1 _11991_ (
    .A1(_00052_),
    .A2(_00516_),
    .B1(addr_i_3_),
    .B2(addr_i_2_),
    .Y(_01671_)
  );
  sg13g2_buf_1 _11992_ (
    .A(_04804_),
    .X(_01672_)
  );
  sg13g2_nand2_1 _11993_ (
    .A(_00117_),
    .B(_00246_),
    .Y(_01673_)
  );
  sg13g2_buf_1 _11994_ (
    .A(_04450_),
    .X(_01674_)
  );
  sg13g2_a22oi_1 _11995_ (
    .A1(_01672_),
    .A2(_01673_),
    .B1(_01674_),
    .B2(addr_i_6_),
    .Y(_01675_)
  );
  sg13g2_nor3_1 _11996_ (
    .A(addr_i_4_),
    .B(_01671_),
    .C(_01675_),
    .Y(_01676_)
  );
  sg13g2_a221oi_1 _11997_ (
    .A1(_06740_),
    .A2(_09226_),
    .B1(_00239_),
    .B2(_09473_),
    .C1(_09271_),
    .Y(_01677_)
  );
  sg13g2_or3_1 _11998_ (
    .A(_00214_),
    .B(_01676_),
    .C(_01677_),
    .X(_01678_)
  );
  sg13g2_o21ai_1 _11999_ (
    .A1(_01665_),
    .A2(_01670_),
    .B1(_01678_),
    .Y(_01679_)
  );
  sg13g2_nand2_1 _12000_ (
    .A(_00511_),
    .B(_01679_),
    .Y(_01681_)
  );
  sg13g2_nand3_1 _12001_ (
    .A(addr_i_11_),
    .B(_01648_),
    .C(_01681_),
    .Y(_01682_)
  );
  sg13g2_nand2_1 _12002_ (
    .A(addr_i_12_),
    .B(_01682_),
    .Y(_01683_)
  );
  sg13g2_nand2_1 _12003_ (
    .A(_09485_),
    .B(_00079_),
    .Y(_01684_)
  );
  sg13g2_a21oi_1 _12004_ (
    .A1(_00427_),
    .A2(_01684_),
    .B1(addr_i_5_),
    .Y(_01685_)
  );
  sg13g2_o21ai_1 _12005_ (
    .A1(_04063_),
    .A2(_00316_),
    .B1(addr_i_3_),
    .Y(_01686_)
  );
  sg13g2_a21o_1 _12006_ (
    .A1(_04285_),
    .A2(_06773_),
    .B1(addr_i_4_),
    .X(_01687_)
  );
  sg13g2_o21ai_1 _12007_ (
    .A1(addr_i_5_),
    .A2(_08100_),
    .B1(_01436_),
    .Y(_01688_)
  );
  sg13g2_nand4_1 _12008_ (
    .A(_01674_),
    .B(_02349_),
    .C(_01687_),
    .D(_01688_),
    .Y(_01689_)
  );
  sg13g2_o21ai_1 _12009_ (
    .A1(_01685_),
    .A2(_01686_),
    .B1(_01689_),
    .Y(_01690_)
  );
  sg13g2_nand2_1 _12010_ (
    .A(_05014_),
    .B(_06530_),
    .Y(_01692_)
  );
  sg13g2_nand3_1 _12011_ (
    .A(addr_i_8_),
    .B(_01690_),
    .C(_01692_),
    .Y(_01693_)
  );
  sg13g2_nand2_1 _12012_ (
    .A(_03380_),
    .B(_07105_),
    .Y(_01694_)
  );
  sg13g2_o21ai_1 _12013_ (
    .A1(_00376_),
    .A2(_00057_),
    .B1(_02514_),
    .Y(_01695_)
  );
  sg13g2_a21oi_1 _12014_ (
    .A1(_01694_),
    .A2(_01695_),
    .B1(addr_i_2_),
    .Y(_01696_)
  );
  sg13g2_xnor2_1 _12015_ (
    .A(addr_i_4_),
    .B(addr_i_6_),
    .Y(_01697_)
  );
  sg13g2_nand3_1 _12016_ (
    .A(_08696_),
    .B(_00316_),
    .C(_07492_),
    .Y(_01698_)
  );
  sg13g2_o21ai_1 _12017_ (
    .A1(_00547_),
    .A2(_00498_),
    .B1(_01698_),
    .Y(_01699_)
  );
  sg13g2_a221oi_1 _12018_ (
    .A1(_01191_),
    .A2(_01697_),
    .B1(_01699_),
    .B2(addr_i_2_),
    .C1(addr_i_8_),
    .Y(_01700_)
  );
  sg13g2_nand2b_1 _12019_ (
    .A_N(_01696_),
    .B(_01700_),
    .Y(_01701_)
  );
  sg13g2_nand2_1 _12020_ (
    .A(_01693_),
    .B(_01701_),
    .Y(_01703_)
  );
  sg13g2_nand2_1 _12021_ (
    .A(_08044_),
    .B(_09485_),
    .Y(_01704_)
  );
  sg13g2_a21oi_1 _12022_ (
    .A1(_09509_),
    .A2(_01704_),
    .B1(_01208_),
    .Y(_01705_)
  );
  sg13g2_nor2_1 _12023_ (
    .A(addr_i_5_),
    .B(_01694_),
    .Y(_01706_)
  );
  sg13g2_a22oi_1 _12024_ (
    .A1(_01231_),
    .A2(_01302_),
    .B1(_01705_),
    .B2(_01706_),
    .Y(_01707_)
  );
  sg13g2_nand2_1 _12025_ (
    .A(_03665_),
    .B(_00676_),
    .Y(_01708_)
  );
  sg13g2_nand2_1 _12026_ (
    .A(addr_i_3_),
    .B(_07658_),
    .Y(_01709_)
  );
  sg13g2_nand3_1 _12027_ (
    .A(_01050_),
    .B(_01708_),
    .C(_01709_),
    .Y(_01710_)
  );
  sg13g2_nor2_1 _12028_ (
    .A(addr_i_7_),
    .B(_02185_),
    .Y(_01711_)
  );
  sg13g2_a221oi_1 _12029_ (
    .A1(addr_i_7_),
    .A2(_01710_),
    .B1(_01711_),
    .B2(_00412_),
    .C1(_07282_),
    .Y(_01712_)
  );
  sg13g2_o21ai_1 _12030_ (
    .A1(addr_i_2_),
    .A2(_01707_),
    .B1(_01712_),
    .Y(_01714_)
  );
  sg13g2_nand2_1 _12031_ (
    .A(_00231_),
    .B(_07956_),
    .Y(_01715_)
  );
  sg13g2_nand2_1 _12032_ (
    .A(_04715_),
    .B(_01715_),
    .Y(_01716_)
  );
  sg13g2_a21oi_1 _12033_ (
    .A1(addr_i_3_),
    .A2(_01716_),
    .B1(_05932_),
    .Y(_01717_)
  );
  sg13g2_nor2_1 _12034_ (
    .A(addr_i_6_),
    .B(_00624_),
    .Y(_01718_)
  );
  sg13g2_o21ai_1 _12035_ (
    .A1(_04284_),
    .A2(_00011_),
    .B1(_01888_),
    .Y(_01719_)
  );
  sg13g2_o21ai_1 _12036_ (
    .A1(_00549_),
    .A2(_01718_),
    .B1(_01719_),
    .Y(_01720_)
  );
  sg13g2_a22oi_1 _12037_ (
    .A1(_00565_),
    .A2(_01720_),
    .B1(_08310_),
    .B2(addr_i_8_),
    .Y(_01721_)
  );
  sg13g2_o21ai_1 _12038_ (
    .A1(addr_i_7_),
    .A2(_01717_),
    .B1(_01721_),
    .Y(_01722_)
  );
  sg13g2_nand3_1 _12039_ (
    .A(addr_i_9_),
    .B(_01714_),
    .C(_01722_),
    .Y(_01723_)
  );
  sg13g2_o21ai_1 _12040_ (
    .A1(addr_i_9_),
    .A2(_01703_),
    .B1(_01723_),
    .Y(_01725_)
  );
  sg13g2_nor3_1 _12041_ (
    .A(addr_i_4_),
    .B(_01867_),
    .C(_09226_),
    .Y(_01726_)
  );
  sg13g2_o21ai_1 _12042_ (
    .A1(_01232_),
    .A2(_01726_),
    .B1(_00067_),
    .Y(_01727_)
  );
  sg13g2_o21ai_1 _12043_ (
    .A1(_01520_),
    .A2(_07050_),
    .B1(_01727_),
    .Y(_01728_)
  );
  sg13g2_nand2_1 _12044_ (
    .A(addr_i_2_),
    .B(_05424_),
    .Y(_01729_)
  );
  sg13g2_nand2_1 _12045_ (
    .A(_00020_),
    .B(_01729_),
    .Y(_01730_)
  );
  sg13g2_a21oi_1 _12046_ (
    .A1(_03919_),
    .A2(_01588_),
    .B1(_03953_),
    .Y(_01731_)
  );
  sg13g2_nor2_1 _12047_ (
    .A(_01592_),
    .B(_04418_),
    .Y(_01732_)
  );
  sg13g2_a22oi_1 _12048_ (
    .A1(addr_i_4_),
    .A2(_01730_),
    .B1(_01731_),
    .B2(_01732_),
    .Y(_01733_)
  );
  sg13g2_nand2_1 _12049_ (
    .A(_07757_),
    .B(_09485_),
    .Y(_01734_)
  );
  sg13g2_o21ai_1 _12050_ (
    .A1(addr_i_3_),
    .A2(_01733_),
    .B1(_01734_),
    .Y(_01736_)
  );
  sg13g2_a22oi_1 _12051_ (
    .A1(addr_i_3_),
    .A2(_01728_),
    .B1(_01736_),
    .B2(_01151_),
    .Y(_01737_)
  );
  sg13g2_buf_1 _12052_ (
    .A(_03413_),
    .X(_01738_)
  );
  sg13g2_a21oi_1 _12053_ (
    .A1(addr_i_5_),
    .A2(_01738_),
    .B1(_00354_),
    .Y(_01739_)
  );
  sg13g2_nand2_1 _12054_ (
    .A(_05169_),
    .B(_00252_),
    .Y(_01740_)
  );
  sg13g2_nand2_1 _12055_ (
    .A(_00927_),
    .B(_01740_),
    .Y(_01741_)
  );
  sg13g2_o21ai_1 _12056_ (
    .A1(_01739_),
    .A2(_01741_),
    .B1(addr_i_6_),
    .Y(_01742_)
  );
  sg13g2_o21ai_1 _12057_ (
    .A1(_00317_),
    .A2(_05557_),
    .B1(_01742_),
    .Y(_01743_)
  );
  sg13g2_nand2b_1 _12058_ (
    .A_N(_01291_),
    .B(_01386_),
    .Y(_01744_)
  );
  sg13g2_nor2_1 _12059_ (
    .A(addr_i_3_),
    .B(addr_i_7_),
    .Y(_01745_)
  );
  sg13g2_buf_1 _12060_ (
    .A(_01745_),
    .X(_01747_)
  );
  sg13g2_a221oi_1 _12061_ (
    .A1(addr_i_3_),
    .A2(_01743_),
    .B1(_01744_),
    .B2(_01747_),
    .C1(addr_i_8_),
    .Y(_01748_)
  );
  sg13g2_nand2_1 _12062_ (
    .A(_08741_),
    .B(_05457_),
    .Y(_01749_)
  );
  sg13g2_nor2_1 _12063_ (
    .A(_00972_),
    .B(_01749_),
    .Y(_01750_)
  );
  sg13g2_a21oi_1 _12064_ (
    .A1(_01047_),
    .A2(_01750_),
    .B1(_00396_),
    .Y(_01751_)
  );
  sg13g2_o21ai_1 _12065_ (
    .A1(_01737_),
    .A2(_01748_),
    .B1(_01751_),
    .Y(_01752_)
  );
  sg13g2_a21oi_1 _12066_ (
    .A1(addr_i_3_),
    .A2(_01254_),
    .B1(_01031_),
    .Y(_01753_)
  );
  sg13g2_nor2_1 _12067_ (
    .A(addr_i_4_),
    .B(_04749_),
    .Y(_01754_)
  );
  sg13g2_a21oi_1 _12068_ (
    .A1(_00565_),
    .A2(_01754_),
    .B1(_01097_),
    .Y(_01755_)
  );
  sg13g2_a21oi_1 _12069_ (
    .A1(addr_i_5_),
    .A2(_01753_),
    .B1(_01755_),
    .Y(_01756_)
  );
  sg13g2_nor2_1 _12070_ (
    .A(addr_i_5_),
    .B(_00770_),
    .Y(_01758_)
  );
  sg13g2_nor2_1 _12071_ (
    .A(_00293_),
    .B(_02536_),
    .Y(_01759_)
  );
  sg13g2_nor4_1 _12072_ (
    .A(_01302_),
    .B(_01758_),
    .C(_01759_),
    .D(_01663_),
    .Y(_01760_)
  );
  sg13g2_a22oi_1 _12073_ (
    .A1(_00610_),
    .A2(_01756_),
    .B1(_01760_),
    .B2(addr_i_9_),
    .Y(_01761_)
  );
  sg13g2_a21oi_1 _12074_ (
    .A1(_01070_),
    .A2(_00453_),
    .B1(_00573_),
    .Y(_01762_)
  );
  sg13g2_a21oi_1 _12075_ (
    .A1(_00386_),
    .A2(_01730_),
    .B1(_01762_),
    .Y(_01763_)
  );
  sg13g2_nor2_1 _12076_ (
    .A(addr_i_3_),
    .B(_01763_),
    .Y(_01764_)
  );
  sg13g2_o21ai_1 _12077_ (
    .A1(addr_i_4_),
    .A2(addr_i_5_),
    .B1(addr_i_6_),
    .Y(_01765_)
  );
  sg13g2_a21oi_1 _12078_ (
    .A1(_00594_),
    .A2(_01765_),
    .B1(_01387_),
    .Y(_01766_)
  );
  sg13g2_nand2_1 _12079_ (
    .A(_00239_),
    .B(_09507_),
    .Y(_01767_)
  );
  sg13g2_o21ai_1 _12080_ (
    .A1(addr_i_7_),
    .A2(_01766_),
    .B1(_01767_),
    .Y(_01769_)
  );
  sg13g2_o21ai_1 _12081_ (
    .A1(_01764_),
    .A2(_01769_),
    .B1(addr_i_8_),
    .Y(_01770_)
  );
  sg13g2_a21oi_1 _12082_ (
    .A1(_01761_),
    .A2(_01770_),
    .B1(addr_i_10_),
    .Y(_01771_)
  );
  sg13g2_a221oi_1 _12083_ (
    .A1(addr_i_10_),
    .A2(_01725_),
    .B1(_01752_),
    .B2(_01771_),
    .C1(addr_i_11_),
    .Y(_01772_)
  );
  sg13g2_buf_1 _12084_ (
    .A(_03731_),
    .X(_01773_)
  );
  sg13g2_buf_1 _12085_ (
    .A(_01773_),
    .X(_01774_)
  );
  sg13g2_o21ai_1 _12086_ (
    .A1(_09094_),
    .A2(_01031_),
    .B1(addr_i_3_),
    .Y(_01775_)
  );
  sg13g2_a21oi_1 _12087_ (
    .A1(_00284_),
    .A2(_00671_),
    .B1(addr_i_3_),
    .Y(_01776_)
  );
  sg13g2_nor2_1 _12088_ (
    .A(_00535_),
    .B(_03314_),
    .Y(_01777_)
  );
  sg13g2_o21ai_1 _12089_ (
    .A1(_01776_),
    .A2(_01777_),
    .B1(addr_i_5_),
    .Y(_01778_)
  );
  sg13g2_nand4_1 _12090_ (
    .A(addr_i_7_),
    .B(_02898_),
    .C(_01775_),
    .D(_01778_),
    .Y(_01780_)
  );
  sg13g2_nand2_1 _12091_ (
    .A(addr_i_8_),
    .B(_01780_),
    .Y(_01781_)
  );
  sg13g2_nor2_1 _12092_ (
    .A(addr_i_3_),
    .B(_03952_),
    .Y(_01782_)
  );
  sg13g2_o21ai_1 _12093_ (
    .A1(_00266_),
    .A2(_01782_),
    .B1(_06375_),
    .Y(_01783_)
  );
  sg13g2_a21oi_1 _12094_ (
    .A1(_00394_),
    .A2(_01783_),
    .B1(addr_i_2_),
    .Y(_01784_)
  );
  sg13g2_a22oi_1 _12095_ (
    .A1(_00743_),
    .A2(_01240_),
    .B1(_01784_),
    .B2(addr_i_7_),
    .Y(_01785_)
  );
  sg13g2_nand3_1 _12096_ (
    .A(_00535_),
    .B(addr_i_6_),
    .C(_00380_),
    .Y(_01786_)
  );
  sg13g2_nor2_1 _12097_ (
    .A(_05856_),
    .B(_05689_),
    .Y(_01787_)
  );
  sg13g2_nor2_1 _12098_ (
    .A(addr_i_7_),
    .B(_01787_),
    .Y(_01788_)
  );
  sg13g2_nand2_1 _12099_ (
    .A(_00581_),
    .B(_01066_),
    .Y(_01789_)
  );
  sg13g2_buf_1 _12100_ (
    .A(_01337_),
    .X(_01791_)
  );
  sg13g2_nand2_1 _12101_ (
    .A(_07282_),
    .B(_01791_),
    .Y(_01792_)
  );
  sg13g2_a221oi_1 _12102_ (
    .A1(_01786_),
    .A2(_01788_),
    .B1(_01789_),
    .B2(_01227_),
    .C1(_01792_),
    .Y(_01793_)
  );
  sg13g2_buf_1 _12103_ (
    .A(_01114_),
    .X(_01794_)
  );
  sg13g2_nand2_1 _12104_ (
    .A(_00593_),
    .B(_00038_),
    .Y(_01795_)
  );
  sg13g2_nand3_1 _12105_ (
    .A(_00414_),
    .B(_00894_),
    .C(_01795_),
    .Y(_01796_)
  );
  sg13g2_nand2_1 _12106_ (
    .A(_01794_),
    .B(_01796_),
    .Y(_01797_)
  );
  sg13g2_a21oi_1 _12107_ (
    .A1(_01793_),
    .A2(_01797_),
    .B1(addr_i_9_),
    .Y(_01798_)
  );
  sg13g2_o21ai_1 _12108_ (
    .A1(_01781_),
    .A2(_01785_),
    .B1(_01798_),
    .Y(_01799_)
  );
  sg13g2_o21ai_1 _12109_ (
    .A1(_03842_),
    .A2(_01954_),
    .B1(_06607_),
    .Y(_01800_)
  );
  sg13g2_o21ai_1 _12110_ (
    .A1(addr_i_3_),
    .A2(_03325_),
    .B1(_01800_),
    .Y(_01802_)
  );
  sg13g2_nor2_1 _12111_ (
    .A(_00030_),
    .B(_00284_),
    .Y(_01803_)
  );
  sg13g2_a22oi_1 _12112_ (
    .A1(addr_i_2_),
    .A2(_01802_),
    .B1(_01803_),
    .B2(addr_i_7_),
    .Y(_01804_)
  );
  sg13g2_a21oi_1 _12113_ (
    .A1(_05745_),
    .A2(_01208_),
    .B1(addr_i_2_),
    .Y(_01805_)
  );
  sg13g2_a22oi_1 _12114_ (
    .A1(addr_i_3_),
    .A2(_01527_),
    .B1(_01459_),
    .B2(addr_i_4_),
    .Y(_01806_)
  );
  sg13g2_o21ai_1 _12115_ (
    .A1(_01805_),
    .A2(_01806_),
    .B1(addr_i_6_),
    .Y(_01807_)
  );
  sg13g2_nand2_1 _12116_ (
    .A(_00956_),
    .B(_00024_),
    .Y(_01808_)
  );
  sg13g2_a22oi_1 _12117_ (
    .A1(_01519_),
    .A2(_01808_),
    .B1(_01660_),
    .B2(_06619_),
    .Y(_01809_)
  );
  sg13g2_nand2_1 _12118_ (
    .A(_01807_),
    .B(_01809_),
    .Y(_01810_)
  );
  sg13g2_nand3b_1 _12119_ (
    .A_N(_01804_),
    .B(addr_i_8_),
    .C(_01810_),
    .Y(_01811_)
  );
  sg13g2_nand2_1 _12120_ (
    .A(addr_i_5_),
    .B(_03314_),
    .Y(_01813_)
  );
  sg13g2_o21ai_1 _12121_ (
    .A1(addr_i_3_),
    .A2(_01628_),
    .B1(_01527_),
    .Y(_01814_)
  );
  sg13g2_buf_1 _12122_ (
    .A(_05678_),
    .X(_01815_)
  );
  sg13g2_a21oi_1 _12123_ (
    .A1(addr_i_6_),
    .A2(_01339_),
    .B1(_01815_),
    .Y(_01816_)
  );
  sg13g2_a221oi_1 _12124_ (
    .A1(_00239_),
    .A2(_01813_),
    .B1(_01814_),
    .B2(addr_i_4_),
    .C1(_01816_),
    .Y(_01817_)
  );
  sg13g2_nand2b_1 _12125_ (
    .A_N(_01817_),
    .B(_00440_),
    .Y(_01818_)
  );
  sg13g2_nor2_1 _12126_ (
    .A(_09510_),
    .B(_00498_),
    .Y(_01819_)
  );
  sg13g2_a21oi_1 _12127_ (
    .A1(_00762_),
    .A2(_00320_),
    .B1(_00151_),
    .Y(_01820_)
  );
  sg13g2_o21ai_1 _12128_ (
    .A1(_01819_),
    .A2(_01820_),
    .B1(_00610_),
    .Y(_01821_)
  );
  sg13g2_nand4_1 _12129_ (
    .A(addr_i_9_),
    .B(_01811_),
    .C(_01818_),
    .D(_01821_),
    .Y(_01822_)
  );
  sg13g2_nand3_1 _12130_ (
    .A(_01774_),
    .B(_01799_),
    .C(_01822_),
    .Y(_01824_)
  );
  sg13g2_nor2_1 _12131_ (
    .A(addr_i_4_),
    .B(_08763_),
    .Y(_01825_)
  );
  sg13g2_nor2_1 _12132_ (
    .A(addr_i_5_),
    .B(_01026_),
    .Y(_01826_)
  );
  sg13g2_o21ai_1 _12133_ (
    .A1(_01825_),
    .A2(_01826_),
    .B1(addr_i_3_),
    .Y(_01827_)
  );
  sg13g2_o21ai_1 _12134_ (
    .A1(_09459_),
    .A2(_00885_),
    .B1(addr_i_2_),
    .Y(_01828_)
  );
  sg13g2_nand2_1 _12135_ (
    .A(_01827_),
    .B(_01828_),
    .Y(_01829_)
  );
  sg13g2_nand2_1 _12136_ (
    .A(_00019_),
    .B(_01834_),
    .Y(_01830_)
  );
  sg13g2_o21ai_1 _12137_ (
    .A1(addr_i_3_),
    .A2(_00079_),
    .B1(_05457_),
    .Y(_01831_)
  );
  sg13g2_a221oi_1 _12138_ (
    .A1(addr_i_3_),
    .A2(_01830_),
    .B1(_01831_),
    .B2(addr_i_5_),
    .C1(addr_i_6_),
    .Y(_01832_)
  );
  sg13g2_a22oi_1 _12139_ (
    .A1(addr_i_6_),
    .A2(_00703_),
    .B1(_01832_),
    .B2(addr_i_7_),
    .Y(_01833_)
  );
  sg13g2_a22oi_1 _12140_ (
    .A1(addr_i_7_),
    .A2(_01829_),
    .B1(_01833_),
    .B2(addr_i_8_),
    .Y(_01835_)
  );
  sg13g2_nor3_1 _12141_ (
    .A(addr_i_3_),
    .B(_08299_),
    .C(_00376_),
    .Y(_01836_)
  );
  sg13g2_buf_1 _12142_ (
    .A(_01292_),
    .X(_01837_)
  );
  sg13g2_a22oi_1 _12143_ (
    .A1(_01528_),
    .A2(_00665_),
    .B1(_01837_),
    .B2(_00822_),
    .Y(_01838_)
  );
  sg13g2_nand2_1 _12144_ (
    .A(addr_i_4_),
    .B(_00329_),
    .Y(_01839_)
  );
  sg13g2_o21ai_1 _12145_ (
    .A1(_01836_),
    .A2(_01838_),
    .B1(_01839_),
    .Y(_01840_)
  );
  sg13g2_nor2_1 _12146_ (
    .A(_07447_),
    .B(_01910_),
    .Y(_01841_)
  );
  sg13g2_o21ai_1 _12147_ (
    .A1(_00324_),
    .A2(_01841_),
    .B1(addr_i_8_),
    .Y(_01842_)
  );
  sg13g2_nand2_1 _12148_ (
    .A(addr_i_3_),
    .B(_01373_),
    .Y(_01843_)
  );
  sg13g2_nand2_1 _12149_ (
    .A(_00697_),
    .B(_01843_),
    .Y(_01844_)
  );
  sg13g2_nor2_1 _12150_ (
    .A(_00030_),
    .B(_04318_),
    .Y(_01846_)
  );
  sg13g2_a22oi_1 _12151_ (
    .A1(_01095_),
    .A2(_01844_),
    .B1(_01846_),
    .B2(_00390_),
    .Y(_01847_)
  );
  sg13g2_a22oi_1 _12152_ (
    .A1(addr_i_7_),
    .A2(_01840_),
    .B1(_01842_),
    .B2(_01847_),
    .Y(_01848_)
  );
  sg13g2_nor2_1 _12153_ (
    .A(_01835_),
    .B(_01848_),
    .Y(_01849_)
  );
  sg13g2_nor2_1 _12154_ (
    .A(_08343_),
    .B(_02733_),
    .Y(_01850_)
  );
  sg13g2_a21oi_1 _12155_ (
    .A1(addr_i_2_),
    .A2(_00819_),
    .B1(_05302_),
    .Y(_01851_)
  );
  sg13g2_o21ai_1 _12156_ (
    .A1(_01850_),
    .A2(_01851_),
    .B1(_04251_),
    .Y(_01852_)
  );
  sg13g2_o21ai_1 _12157_ (
    .A1(_00938_),
    .A2(_00079_),
    .B1(_00020_),
    .Y(_01853_)
  );
  sg13g2_a21oi_1 _12158_ (
    .A1(_05867_),
    .A2(_01853_),
    .B1(_08575_),
    .Y(_01854_)
  );
  sg13g2_a21oi_1 _12159_ (
    .A1(_01852_),
    .A2(_01854_),
    .B1(addr_i_7_),
    .Y(_01855_)
  );
  sg13g2_nand2_1 _12160_ (
    .A(_00072_),
    .B(_00959_),
    .Y(_01857_)
  );
  sg13g2_a21oi_1 _12161_ (
    .A1(_02656_),
    .A2(_01857_),
    .B1(_06895_),
    .Y(_01858_)
  );
  sg13g2_nor2_1 _12162_ (
    .A(_01855_),
    .B(_01858_),
    .Y(_01859_)
  );
  sg13g2_o21ai_1 _12163_ (
    .A1(_00807_),
    .A2(_01859_),
    .B1(addr_i_11_),
    .Y(_01860_)
  );
  sg13g2_buf_1 _12164_ (
    .A(_01310_),
    .X(_01861_)
  );
  sg13g2_o21ai_1 _12165_ (
    .A1(_06154_),
    .A2(_01031_),
    .B1(_05867_),
    .Y(_01862_)
  );
  sg13g2_nor2_1 _12166_ (
    .A(_01976_),
    .B(_02207_),
    .Y(_01863_)
  );
  sg13g2_o21ai_1 _12167_ (
    .A1(_01459_),
    .A2(_01863_),
    .B1(addr_i_4_),
    .Y(_01864_)
  );
  sg13g2_nand3_1 _12168_ (
    .A(_00148_),
    .B(_01862_),
    .C(_01864_),
    .Y(_01865_)
  );
  sg13g2_a21oi_1 _12169_ (
    .A1(_08930_),
    .A2(_02887_),
    .B1(addr_i_3_),
    .Y(_01866_)
  );
  sg13g2_a21oi_1 _12170_ (
    .A1(addr_i_3_),
    .A2(_03325_),
    .B1(_01866_),
    .Y(_01868_)
  );
  sg13g2_nor2_1 _12171_ (
    .A(addr_i_4_),
    .B(_00663_),
    .Y(_01869_)
  );
  sg13g2_o21ai_1 _12172_ (
    .A1(_01024_),
    .A2(_01869_),
    .B1(addr_i_3_),
    .Y(_01870_)
  );
  sg13g2_o21ai_1 _12173_ (
    .A1(addr_i_2_),
    .A2(_01868_),
    .B1(_01870_),
    .Y(_01871_)
  );
  sg13g2_buf_1 _12174_ (
    .A(_00287_),
    .X(_01872_)
  );
  sg13g2_nand3_1 _12175_ (
    .A(addr_i_4_),
    .B(_01872_),
    .C(_01795_),
    .Y(_01873_)
  );
  sg13g2_a21oi_1 _12176_ (
    .A1(_00762_),
    .A2(_01873_),
    .B1(_04672_),
    .Y(_01874_)
  );
  sg13g2_a221oi_1 _12177_ (
    .A1(_01861_),
    .A2(_01865_),
    .B1(_01871_),
    .B2(_00708_),
    .C1(_01874_),
    .Y(_01875_)
  );
  sg13g2_nor2_1 _12178_ (
    .A(_01211_),
    .B(_01875_),
    .Y(_01876_)
  );
  sg13g2_a22oi_1 _12179_ (
    .A1(_05214_),
    .A2(_01849_),
    .B1(_01860_),
    .B2(_01876_),
    .Y(_01877_)
  );
  sg13g2_a21oi_1 _12180_ (
    .A1(_01824_),
    .A2(_01877_),
    .B1(addr_i_12_),
    .Y(_01879_)
  );
  sg13g2_nand2b_1 _12181_ (
    .A_N(_01772_),
    .B(_01879_),
    .Y(_01880_)
  );
  sg13g2_o21ai_1 _12182_ (
    .A1(_01642_),
    .A2(_01683_),
    .B1(_01880_),
    .Y(data_o_13_)
  );
  sg13g2_buf_1 _12183_ (
    .A(_03380_),
    .X(_01881_)
  );
  sg13g2_nor2_1 _12184_ (
    .A(_01881_),
    .B(_01456_),
    .Y(_01882_)
  );
  sg13g2_o21ai_1 _12185_ (
    .A1(_01302_),
    .A2(_01179_),
    .B1(_01882_),
    .Y(_01883_)
  );
  sg13g2_a21oi_1 _12186_ (
    .A1(_00529_),
    .A2(_01883_),
    .B1(addr_i_8_),
    .Y(_01884_)
  );
  sg13g2_a221oi_1 _12187_ (
    .A1(_00238_),
    .A2(_00665_),
    .B1(_01244_),
    .B2(_00687_),
    .C1(_06264_),
    .Y(_01885_)
  );
  sg13g2_nand2_1 _12188_ (
    .A(addr_i_6_),
    .B(_02218_),
    .Y(_01886_)
  );
  sg13g2_a22oi_1 _12189_ (
    .A1(addr_i_2_),
    .A2(_01886_),
    .B1(_00746_),
    .B2(addr_i_4_),
    .Y(_01887_)
  );
  sg13g2_a22oi_1 _12190_ (
    .A1(addr_i_4_),
    .A2(_01885_),
    .B1(_01887_),
    .B2(addr_i_7_),
    .Y(_01889_)
  );
  sg13g2_a21oi_1 _12191_ (
    .A1(_06508_),
    .A2(_01465_),
    .B1(_00053_),
    .Y(_01890_)
  );
  sg13g2_nor2_1 _12192_ (
    .A(_01889_),
    .B(_01890_),
    .Y(_01891_)
  );
  sg13g2_buf_1 _12193_ (
    .A(_00262_),
    .X(_01892_)
  );
  sg13g2_o21ai_1 _12194_ (
    .A1(addr_i_2_),
    .A2(_03853_),
    .B1(_00822_),
    .Y(_01893_)
  );
  sg13g2_o21ai_1 _12195_ (
    .A1(addr_i_5_),
    .A2(_00238_),
    .B1(addr_i_4_),
    .Y(_01894_)
  );
  sg13g2_nand3_1 _12196_ (
    .A(_09476_),
    .B(_01893_),
    .C(_01894_),
    .Y(_01895_)
  );
  sg13g2_nor2_1 _12197_ (
    .A(addr_i_3_),
    .B(_01373_),
    .Y(_01896_)
  );
  sg13g2_o21ai_1 _12198_ (
    .A1(_05258_),
    .A2(_01896_),
    .B1(addr_i_4_),
    .Y(_01897_)
  );
  sg13g2_a21o_1 _12199_ (
    .A1(_00762_),
    .A2(_01795_),
    .B1(addr_i_4_),
    .X(_01898_)
  );
  sg13g2_a21oi_1 _12200_ (
    .A1(_01897_),
    .A2(_01898_),
    .B1(_01481_),
    .Y(_01900_)
  );
  sg13g2_nor2_1 _12201_ (
    .A(addr_i_2_),
    .B(_08166_),
    .Y(_01901_)
  );
  sg13g2_nor2_1 _12202_ (
    .A(addr_i_3_),
    .B(_02602_),
    .Y(_01902_)
  );
  sg13g2_a22oi_1 _12203_ (
    .A1(addr_i_3_),
    .A2(_01901_),
    .B1(_01902_),
    .B2(_00617_),
    .Y(_01903_)
  );
  sg13g2_a21oi_1 _12204_ (
    .A1(_00381_),
    .A2(_02470_),
    .B1(_00052_),
    .Y(_01904_)
  );
  sg13g2_nor2_1 _12205_ (
    .A(_05888_),
    .B(_01904_),
    .Y(_01905_)
  );
  sg13g2_o21ai_1 _12206_ (
    .A1(_00230_),
    .A2(_01903_),
    .B1(_01905_),
    .Y(_01906_)
  );
  sg13g2_a22oi_1 _12207_ (
    .A1(_01892_),
    .A2(_01895_),
    .B1(_01900_),
    .B2(_01906_),
    .Y(_01907_)
  );
  sg13g2_a21oi_1 _12208_ (
    .A1(_01884_),
    .A2(_01891_),
    .B1(_01907_),
    .Y(_01908_)
  );
  sg13g2_xnor2_1 _12209_ (
    .A(_01548_),
    .B(_01901_),
    .Y(_01909_)
  );
  sg13g2_nand2_1 _12210_ (
    .A(addr_i_4_),
    .B(addr_i_8_),
    .Y(_01911_)
  );
  sg13g2_buf_1 _12211_ (
    .A(_01084_),
    .X(_01912_)
  );
  sg13g2_o21ai_1 _12212_ (
    .A1(_00150_),
    .A2(_01911_),
    .B1(_01912_),
    .Y(_01913_)
  );
  sg13g2_nand2b_1 _12213_ (
    .A_N(addr_i_4_),
    .B(addr_i_8_),
    .Y(_01914_)
  );
  sg13g2_nor2_1 _12214_ (
    .A(_00329_),
    .B(_01914_),
    .Y(_01915_)
  );
  sg13g2_a22oi_1 _12215_ (
    .A1(addr_i_6_),
    .A2(_01909_),
    .B1(_01913_),
    .B2(_01915_),
    .Y(_01916_)
  );
  sg13g2_nor2_1 _12216_ (
    .A(addr_i_8_),
    .B(addr_i_6_),
    .Y(_01917_)
  );
  sg13g2_nand2_1 _12217_ (
    .A(_01215_),
    .B(_01917_),
    .Y(_01918_)
  );
  sg13g2_nand2_1 _12218_ (
    .A(_01367_),
    .B(_01918_),
    .Y(_01919_)
  );
  sg13g2_nor2b_1 _12219_ (
    .A(addr_i_6_),
    .B_N(addr_i_8_),
    .Y(_01920_)
  );
  sg13g2_o21ai_1 _12220_ (
    .A1(_08896_),
    .A2(_01588_),
    .B1(_01589_),
    .Y(_01922_)
  );
  sg13g2_nor2_1 _12221_ (
    .A(addr_i_8_),
    .B(_03446_),
    .Y(_01923_)
  );
  sg13g2_a22oi_1 _12222_ (
    .A1(_06220_),
    .A2(_01920_),
    .B1(_01922_),
    .B2(_01923_),
    .Y(_01924_)
  );
  sg13g2_nor2_1 _12223_ (
    .A(_00910_),
    .B(_01924_),
    .Y(_01925_)
  );
  sg13g2_a21oi_1 _12224_ (
    .A1(addr_i_5_),
    .A2(_01919_),
    .B1(_01925_),
    .Y(_01926_)
  );
  sg13g2_o21ai_1 _12225_ (
    .A1(addr_i_3_),
    .A2(_01916_),
    .B1(_01926_),
    .Y(_01927_)
  );
  sg13g2_or2_1 _12226_ (
    .A(addr_i_8_),
    .B(addr_i_6_),
    .X(_01928_)
  );
  sg13g2_nor2_1 _12227_ (
    .A(_00744_),
    .B(_01928_),
    .Y(_01929_)
  );
  sg13g2_o21ai_1 _12228_ (
    .A1(_06021_),
    .A2(_01929_),
    .B1(_00594_),
    .Y(_01930_)
  );
  sg13g2_nand2_1 _12229_ (
    .A(_01918_),
    .B(_01930_),
    .Y(_01931_)
  );
  sg13g2_nand2b_1 _12230_ (
    .A_N(addr_i_6_),
    .B(addr_i_8_),
    .Y(_01933_)
  );
  sg13g2_o21ai_1 _12231_ (
    .A1(_00224_),
    .A2(_01933_),
    .B1(addr_i_7_),
    .Y(_01934_)
  );
  sg13g2_buf_1 _12232_ (
    .A(_09491_),
    .X(_01935_)
  );
  sg13g2_nor2b_1 _12233_ (
    .A(addr_i_8_),
    .B_N(addr_i_6_),
    .Y(_01936_)
  );
  sg13g2_nand2_1 _12234_ (
    .A(addr_i_2_),
    .B(_01936_),
    .Y(_01937_)
  );
  sg13g2_a21o_1 _12235_ (
    .A1(_01933_),
    .A2(_01937_),
    .B1(_08155_),
    .X(_01938_)
  );
  sg13g2_a221oi_1 _12236_ (
    .A1(_01528_),
    .A2(_01920_),
    .B1(_01936_),
    .B2(_01308_),
    .C1(_00485_),
    .Y(_01939_)
  );
  sg13g2_a22oi_1 _12237_ (
    .A1(_01935_),
    .A2(_01938_),
    .B1(_01939_),
    .B2(addr_i_5_),
    .Y(_01940_)
  );
  sg13g2_a22oi_1 _12238_ (
    .A1(addr_i_5_),
    .A2(_01931_),
    .B1(_01934_),
    .B2(_01940_),
    .Y(_01941_)
  );
  sg13g2_a22oi_1 _12239_ (
    .A1(_05834_),
    .A2(_01927_),
    .B1(_01941_),
    .B2(addr_i_9_),
    .Y(_01942_)
  );
  sg13g2_a22oi_1 _12240_ (
    .A1(addr_i_9_),
    .A2(_01908_),
    .B1(_01942_),
    .B2(addr_i_10_),
    .Y(_01944_)
  );
  sg13g2_nand2_1 _12241_ (
    .A(_04119_),
    .B(_04284_),
    .Y(_01945_)
  );
  sg13g2_nand2_1 _12242_ (
    .A(addr_i_3_),
    .B(_05225_),
    .Y(_01946_)
  );
  sg13g2_nand2_1 _12243_ (
    .A(_01945_),
    .B(_01946_),
    .Y(_01947_)
  );
  sg13g2_nand2_1 _12244_ (
    .A(_00064_),
    .B(_01680_),
    .Y(_01948_)
  );
  sg13g2_nand2_1 _12245_ (
    .A(_04904_),
    .B(_06485_),
    .Y(_01949_)
  );
  sg13g2_nand2_1 _12246_ (
    .A(addr_i_2_),
    .B(_01949_),
    .Y(_01950_)
  );
  sg13g2_nand3_1 _12247_ (
    .A(_00520_),
    .B(_01948_),
    .C(_01950_),
    .Y(_01951_)
  );
  sg13g2_o21ai_1 _12248_ (
    .A1(_01160_),
    .A2(_01791_),
    .B1(addr_i_8_),
    .Y(_01952_)
  );
  sg13g2_a221oi_1 _12249_ (
    .A1(addr_i_5_),
    .A2(_01947_),
    .B1(_01951_),
    .B2(_00157_),
    .C1(_01952_),
    .Y(_01953_)
  );
  sg13g2_nand2_1 _12250_ (
    .A(_01603_),
    .B(_00433_),
    .Y(_01955_)
  );
  sg13g2_a21oi_1 _12251_ (
    .A1(_00316_),
    .A2(_02459_),
    .B1(addr_i_5_),
    .Y(_01956_)
  );
  sg13g2_nor2_1 _12252_ (
    .A(_01976_),
    .B(_00819_),
    .Y(_01957_)
  );
  sg13g2_a22oi_1 _12253_ (
    .A1(addr_i_3_),
    .A2(_01955_),
    .B1(_01956_),
    .B2(_01957_),
    .Y(_01958_)
  );
  sg13g2_nand2b_1 _12254_ (
    .A_N(_01958_),
    .B(addr_i_4_),
    .Y(_01959_)
  );
  sg13g2_o21ai_1 _12255_ (
    .A1(addr_i_6_),
    .A2(addr_i_5_),
    .B1(addr_i_3_),
    .Y(_01960_)
  );
  sg13g2_a22oi_1 _12256_ (
    .A1(_01368_),
    .A2(_01960_),
    .B1(_00122_),
    .B2(_00930_),
    .Y(_01961_)
  );
  sg13g2_nor2_1 _12257_ (
    .A(_07160_),
    .B(_00718_),
    .Y(_01962_)
  );
  sg13g2_a221oi_1 _12258_ (
    .A1(_09127_),
    .A2(_00400_),
    .B1(_00442_),
    .B2(_00001_),
    .C1(_01962_),
    .Y(_01963_)
  );
  sg13g2_nor2b_1 _12259_ (
    .A(_01961_),
    .B_N(_01963_),
    .Y(_01964_)
  );
  sg13g2_nor2_1 _12260_ (
    .A(addr_i_7_),
    .B(_06530_),
    .Y(_01966_)
  );
  sg13g2_nand2_1 _12261_ (
    .A(addr_i_4_),
    .B(_01856_),
    .Y(_01967_)
  );
  sg13g2_o21ai_1 _12262_ (
    .A1(addr_i_4_),
    .A2(_01966_),
    .B1(_01967_),
    .Y(_01968_)
  );
  sg13g2_nand2_1 _12263_ (
    .A(addr_i_3_),
    .B(_01968_),
    .Y(_01969_)
  );
  sg13g2_buf_1 _12264_ (
    .A(_08156_),
    .X(_01970_)
  );
  sg13g2_nand2_1 _12265_ (
    .A(_01065_),
    .B(_02887_),
    .Y(_01971_)
  );
  sg13g2_buf_1 _12266_ (
    .A(_00624_),
    .X(_01972_)
  );
  sg13g2_a22oi_1 _12267_ (
    .A1(_01970_),
    .A2(_01971_),
    .B1(_01972_),
    .B2(addr_i_2_),
    .Y(_01973_)
  );
  sg13g2_a21oi_1 _12268_ (
    .A1(_01969_),
    .A2(_01973_),
    .B1(addr_i_8_),
    .Y(_01974_)
  );
  sg13g2_a221oi_1 _12269_ (
    .A1(_01953_),
    .A2(_01959_),
    .B1(_01964_),
    .B2(_01974_),
    .C1(addr_i_9_),
    .Y(_01975_)
  );
  sg13g2_nor2_1 _12270_ (
    .A(_02371_),
    .B(_06851_),
    .Y(_01977_)
  );
  sg13g2_a21oi_1 _12271_ (
    .A1(_04318_),
    .A2(_00246_),
    .B1(_04362_),
    .Y(_01978_)
  );
  sg13g2_o21ai_1 _12272_ (
    .A1(_01977_),
    .A2(_01978_),
    .B1(addr_i_3_),
    .Y(_01979_)
  );
  sg13g2_o21ai_1 _12273_ (
    .A1(_00246_),
    .A2(_02591_),
    .B1(_00016_),
    .Y(_01980_)
  );
  sg13g2_a21oi_1 _12274_ (
    .A1(_00483_),
    .A2(_01980_),
    .B1(_06939_),
    .Y(_01981_)
  );
  sg13g2_a21oi_1 _12275_ (
    .A1(_01979_),
    .A2(_01981_),
    .B1(addr_i_6_),
    .Y(_01982_)
  );
  sg13g2_nand2_1 _12276_ (
    .A(addr_i_4_),
    .B(_01055_),
    .Y(_01983_)
  );
  sg13g2_a21o_1 _12277_ (
    .A1(_00249_),
    .A2(_01983_),
    .B1(addr_i_5_),
    .X(_01984_)
  );
  sg13g2_a21oi_1 _12278_ (
    .A1(_01691_),
    .A2(_01984_),
    .B1(addr_i_3_),
    .Y(_01985_)
  );
  sg13g2_nor2_1 _12279_ (
    .A(_09038_),
    .B(_00462_),
    .Y(_01986_)
  );
  sg13g2_o21ai_1 _12280_ (
    .A1(_01507_),
    .A2(_01986_),
    .B1(addr_i_4_),
    .Y(_01988_)
  );
  sg13g2_nand2_1 _12281_ (
    .A(_00112_),
    .B(_01988_),
    .Y(_01989_)
  );
  sg13g2_o21ai_1 _12282_ (
    .A1(addr_i_2_),
    .A2(_00624_),
    .B1(_00679_),
    .Y(_01990_)
  );
  sg13g2_a21oi_1 _12283_ (
    .A1(addr_i_3_),
    .A2(_01990_),
    .B1(_01127_),
    .Y(_01991_)
  );
  sg13g2_nor2_1 _12284_ (
    .A(_04251_),
    .B(_01991_),
    .Y(_01992_)
  );
  sg13g2_nor4_1 _12285_ (
    .A(_01982_),
    .B(_01985_),
    .C(_01989_),
    .D(_01992_),
    .Y(_01993_)
  );
  sg13g2_a21oi_1 _12286_ (
    .A1(_06496_),
    .A2(_06972_),
    .B1(_04450_),
    .Y(_01994_)
  );
  sg13g2_a21oi_1 _12287_ (
    .A1(_02053_),
    .A2(_03743_),
    .B1(_00117_),
    .Y(_01995_)
  );
  sg13g2_o21ai_1 _12288_ (
    .A1(_01994_),
    .A2(_01995_),
    .B1(addr_i_2_),
    .Y(_01996_)
  );
  sg13g2_nand3_1 _12289_ (
    .A(_01331_),
    .B(_09149_),
    .C(_01996_),
    .Y(_01997_)
  );
  sg13g2_o21ai_1 _12290_ (
    .A1(_03139_),
    .A2(_04782_),
    .B1(addr_i_3_),
    .Y(_01999_)
  );
  sg13g2_nand4_1 _12291_ (
    .A(addr_i_8_),
    .B(_01791_),
    .C(_00928_),
    .D(_01999_),
    .Y(_02000_)
  );
  sg13g2_nand2_1 _12292_ (
    .A(addr_i_3_),
    .B(_00879_),
    .Y(_02001_)
  );
  sg13g2_nand2_1 _12293_ (
    .A(_01153_),
    .B(_07492_),
    .Y(_02002_)
  );
  sg13g2_a21oi_1 _12294_ (
    .A1(_02001_),
    .A2(_02002_),
    .B1(addr_i_7_),
    .Y(_02003_)
  );
  sg13g2_a22oi_1 _12295_ (
    .A1(addr_i_4_),
    .A2(_01997_),
    .B1(_02000_),
    .B2(_02003_),
    .Y(_02004_)
  );
  sg13g2_o21ai_1 _12296_ (
    .A1(_01993_),
    .A2(_02004_),
    .B1(addr_i_9_),
    .Y(_02005_)
  );
  sg13g2_nand3b_1 _12297_ (
    .A_N(_01975_),
    .B(addr_i_10_),
    .C(_02005_),
    .Y(_02006_)
  );
  sg13g2_nand2_1 _12298_ (
    .A(_01640_),
    .B(_02006_),
    .Y(_02007_)
  );
  sg13g2_nor2_1 _12299_ (
    .A(addr_i_2_),
    .B(_00665_),
    .Y(_02008_)
  );
  sg13g2_nor2_1 _12300_ (
    .A(_06851_),
    .B(_08796_),
    .Y(_02010_)
  );
  sg13g2_o21ai_1 _12301_ (
    .A1(_02008_),
    .A2(_02010_),
    .B1(_00116_),
    .Y(_02011_)
  );
  sg13g2_buf_1 _12302_ (
    .A(_00413_),
    .X(_02012_)
  );
  sg13g2_nand3_1 _12303_ (
    .A(_02012_),
    .B(_07790_),
    .C(_01872_),
    .Y(_02013_)
  );
  sg13g2_nor3_1 _12304_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .C(_00550_),
    .Y(_02014_)
  );
  sg13g2_nor2_1 _12305_ (
    .A(addr_i_3_),
    .B(_03842_),
    .Y(_02015_)
  );
  sg13g2_o21ai_1 _12306_ (
    .A1(_00155_),
    .A2(_02015_),
    .B1(_07934_),
    .Y(_02016_)
  );
  sg13g2_a221oi_1 _12307_ (
    .A1(addr_i_4_),
    .A2(_02013_),
    .B1(_02014_),
    .B2(addr_i_3_),
    .C1(_02016_),
    .Y(_02017_)
  );
  sg13g2_nor2_1 _12308_ (
    .A(_00009_),
    .B(_00494_),
    .Y(_02018_)
  );
  sg13g2_xnor2_1 _12309_ (
    .A(addr_i_2_),
    .B(_02018_),
    .Y(_02019_)
  );
  sg13g2_nand2_1 _12310_ (
    .A(_00260_),
    .B(_08254_),
    .Y(_02021_)
  );
  sg13g2_a22oi_1 _12311_ (
    .A1(addr_i_4_),
    .A2(_02021_),
    .B1(_07591_),
    .B2(addr_i_6_),
    .Y(_02022_)
  );
  sg13g2_a221oi_1 _12312_ (
    .A1(addr_i_8_),
    .A2(_01580_),
    .B1(_00321_),
    .B2(_02022_),
    .C1(addr_i_9_),
    .Y(_02023_)
  );
  sg13g2_o21ai_1 _12313_ (
    .A1(_01663_),
    .A2(_02019_),
    .B1(_02023_),
    .Y(_02024_)
  );
  sg13g2_nand3_1 _12314_ (
    .A(addr_i_3_),
    .B(_00391_),
    .C(_00039_),
    .Y(_02025_)
  );
  sg13g2_nor2_1 _12315_ (
    .A(_01384_),
    .B(_00521_),
    .Y(_02026_)
  );
  sg13g2_nor2_1 _12316_ (
    .A(addr_i_6_),
    .B(_02026_),
    .Y(_02027_)
  );
  sg13g2_nand2_1 _12317_ (
    .A(_01881_),
    .B(_01104_),
    .Y(_02028_)
  );
  sg13g2_a221oi_1 _12318_ (
    .A1(_02025_),
    .A2(_02027_),
    .B1(_02028_),
    .B2(addr_i_6_),
    .C1(_00802_),
    .Y(_02029_)
  );
  sg13g2_a22oi_1 _12319_ (
    .A1(_02011_),
    .A2(_02017_),
    .B1(_02024_),
    .B2(_02029_),
    .Y(_02030_)
  );
  sg13g2_nand2_1 _12320_ (
    .A(_03908_),
    .B(_00664_),
    .Y(_02032_)
  );
  sg13g2_nand2_1 _12321_ (
    .A(_00846_),
    .B(_02032_),
    .Y(_02033_)
  );
  sg13g2_o21ai_1 _12322_ (
    .A1(addr_i_3_),
    .A2(_00791_),
    .B1(_00789_),
    .Y(_02034_)
  );
  sg13g2_a21o_1 _12323_ (
    .A1(_01310_),
    .A2(_02033_),
    .B1(_02034_),
    .X(_02035_)
  );
  sg13g2_a21oi_1 _12324_ (
    .A1(addr_i_9_),
    .A2(_02035_),
    .B1(addr_i_10_),
    .Y(_02036_)
  );
  sg13g2_nor2b_1 _12325_ (
    .A(_02030_),
    .B_N(_02036_),
    .Y(_02037_)
  );
  sg13g2_o21ai_1 _12326_ (
    .A1(addr_i_3_),
    .A2(_01091_),
    .B1(_01493_),
    .Y(_02038_)
  );
  sg13g2_a21oi_1 _12327_ (
    .A1(_00846_),
    .A2(_02032_),
    .B1(addr_i_7_),
    .Y(_02039_)
  );
  sg13g2_buf_1 _12328_ (
    .A(_00807_),
    .X(_02040_)
  );
  sg13g2_a22oi_1 _12329_ (
    .A1(addr_i_7_),
    .A2(_02038_),
    .B1(_02039_),
    .B2(_02040_),
    .Y(_02041_)
  );
  sg13g2_o21ai_1 _12330_ (
    .A1(_02037_),
    .A2(_02041_),
    .B1(addr_i_11_),
    .Y(_02043_)
  );
  sg13g2_o21ai_1 _12331_ (
    .A1(_01944_),
    .A2(_02007_),
    .B1(_02043_),
    .Y(_02044_)
  );
  sg13g2_o21ai_1 _12332_ (
    .A1(_04063_),
    .A2(_06176_),
    .B1(_01050_),
    .Y(_02045_)
  );
  sg13g2_a221oi_1 _12333_ (
    .A1(_01231_),
    .A2(_01215_),
    .B1(_02045_),
    .B2(addr_i_7_),
    .C1(addr_i_3_),
    .Y(_02046_)
  );
  sg13g2_nand2_1 _12334_ (
    .A(_01153_),
    .B(_03128_),
    .Y(_02047_)
  );
  sg13g2_nand2_1 _12335_ (
    .A(_00303_),
    .B(_00038_),
    .Y(_02048_)
  );
  sg13g2_nand3_1 _12336_ (
    .A(_00863_),
    .B(_02047_),
    .C(_02048_),
    .Y(_02049_)
  );
  sg13g2_a221oi_1 _12337_ (
    .A1(_01159_),
    .A2(_01445_),
    .B1(_02049_),
    .B2(_03820_),
    .C1(_00190_),
    .Y(_02050_)
  );
  sg13g2_or2_1 _12338_ (
    .A(_02046_),
    .B(_02050_),
    .X(_02051_)
  );
  sg13g2_nand2_1 _12339_ (
    .A(_01461_),
    .B(_04860_),
    .Y(_02052_)
  );
  sg13g2_nand3_1 _12340_ (
    .A(_02930_),
    .B(_00368_),
    .C(_02052_),
    .Y(_02054_)
  );
  sg13g2_nor2_1 _12341_ (
    .A(_01055_),
    .B(_01625_),
    .Y(_02055_)
  );
  sg13g2_a22oi_1 _12342_ (
    .A1(addr_i_4_),
    .A2(_00292_),
    .B1(_04506_),
    .B2(_02055_),
    .Y(_02056_)
  );
  sg13g2_nor2_1 _12343_ (
    .A(addr_i_6_),
    .B(_00495_),
    .Y(_02057_)
  );
  sg13g2_a21oi_1 _12344_ (
    .A1(_00211_),
    .A2(_00739_),
    .B1(addr_i_4_),
    .Y(_02058_)
  );
  sg13g2_a221oi_1 _12345_ (
    .A1(_00375_),
    .A2(_01064_),
    .B1(_02057_),
    .B2(_01580_),
    .C1(_02058_),
    .Y(_02059_)
  );
  sg13g2_o21ai_1 _12346_ (
    .A1(addr_i_3_),
    .A2(_02056_),
    .B1(_02059_),
    .Y(_02060_)
  );
  sg13g2_a22oi_1 _12347_ (
    .A1(_00779_),
    .A2(_02054_),
    .B1(_02060_),
    .B2(addr_i_8_),
    .Y(_02061_)
  );
  sg13g2_a21oi_1 _12348_ (
    .A1(addr_i_8_),
    .A2(_02051_),
    .B1(_02061_),
    .Y(_02062_)
  );
  sg13g2_buf_1 _12349_ (
    .A(_06143_),
    .X(_02063_)
  );
  sg13g2_mux2_1 _12350_ (
    .A0(_08089_),
    .A1(_00086_),
    .S(_05845_),
    .X(_02065_)
  );
  sg13g2_nand2_1 _12351_ (
    .A(addr_i_3_),
    .B(_00086_),
    .Y(_02066_)
  );
  sg13g2_o21ai_1 _12352_ (
    .A1(addr_i_6_),
    .A2(_02065_),
    .B1(_02066_),
    .Y(_02067_)
  );
  sg13g2_a21oi_1 _12353_ (
    .A1(_02063_),
    .A2(_02067_),
    .B1(_01627_),
    .Y(_02068_)
  );
  sg13g2_and4_1 _12354_ (
    .A(addr_i_4_),
    .B(addr_i_7_),
    .C(addr_i_6_),
    .D(addr_i_5_),
    .X(_02069_)
  );
  sg13g2_o21ai_1 _12355_ (
    .A1(_07105_),
    .A2(_02069_),
    .B1(addr_i_3_),
    .Y(_02070_)
  );
  sg13g2_o21ai_1 _12356_ (
    .A1(_05745_),
    .A2(_00404_),
    .B1(_02070_),
    .Y(_02071_)
  );
  sg13g2_nor3_1 _12357_ (
    .A(_00692_),
    .B(_00381_),
    .C(_01585_),
    .Y(_02072_)
  );
  sg13g2_a22oi_1 _12358_ (
    .A1(addr_i_2_),
    .A2(_02071_),
    .B1(_02072_),
    .B2(_05888_),
    .Y(_02073_)
  );
  sg13g2_o21ai_1 _12359_ (
    .A1(addr_i_4_),
    .A2(_02068_),
    .B1(_02073_),
    .Y(_02074_)
  );
  sg13g2_buf_1 _12360_ (
    .A(_08453_),
    .X(_02076_)
  );
  sg13g2_nand2_1 _12361_ (
    .A(addr_i_3_),
    .B(_00495_),
    .Y(_02077_)
  );
  sg13g2_a21oi_1 _12362_ (
    .A1(addr_i_7_),
    .A2(_02077_),
    .B1(addr_i_4_),
    .Y(_02078_)
  );
  sg13g2_a22oi_1 _12363_ (
    .A1(_03820_),
    .A2(_02076_),
    .B1(_02078_),
    .B2(_01660_),
    .Y(_02079_)
  );
  sg13g2_nand2_1 _12364_ (
    .A(_03953_),
    .B(_01222_),
    .Y(_02080_)
  );
  sg13g2_nor2_1 _12365_ (
    .A(_08885_),
    .B(_01375_),
    .Y(_02081_)
  );
  sg13g2_nand2_1 _12366_ (
    .A(_04528_),
    .B(_09506_),
    .Y(_02082_)
  );
  sg13g2_o21ai_1 _12367_ (
    .A1(addr_i_7_),
    .A2(_02081_),
    .B1(_02082_),
    .Y(_02083_)
  );
  sg13g2_a221oi_1 _12368_ (
    .A1(_00244_),
    .A2(_02080_),
    .B1(_02083_),
    .B2(_02404_),
    .C1(addr_i_8_),
    .Y(_02084_)
  );
  sg13g2_o21ai_1 _12369_ (
    .A1(addr_i_6_),
    .A2(_02079_),
    .B1(_02084_),
    .Y(_02085_)
  );
  sg13g2_nand2_1 _12370_ (
    .A(_02074_),
    .B(_02085_),
    .Y(_02087_)
  );
  sg13g2_or3_1 _12371_ (
    .A(addr_i_7_),
    .B(addr_i_6_),
    .C(addr_i_5_),
    .X(_02088_)
  );
  sg13g2_buf_1 _12372_ (
    .A(_02088_),
    .X(_02089_)
  );
  sg13g2_nand2_1 _12373_ (
    .A(_02371_),
    .B(_02089_),
    .Y(_02090_)
  );
  sg13g2_nor2_1 _12374_ (
    .A(_06496_),
    .B(_05169_),
    .Y(_02091_)
  );
  sg13g2_nor2_1 _12375_ (
    .A(_05546_),
    .B(_04893_),
    .Y(_02092_)
  );
  sg13g2_a221oi_1 _12376_ (
    .A1(_01888_),
    .A2(_02090_),
    .B1(_02091_),
    .B2(_01215_),
    .C1(_02092_),
    .Y(_02093_)
  );
  sg13g2_nand2_1 _12377_ (
    .A(_09501_),
    .B(_00184_),
    .Y(_02094_)
  );
  sg13g2_nand3_1 _12378_ (
    .A(_06364_),
    .B(addr_i_5_),
    .C(_00406_),
    .Y(_02095_)
  );
  sg13g2_a21oi_1 _12379_ (
    .A1(_02094_),
    .A2(_02095_),
    .B1(addr_i_3_),
    .Y(_02096_)
  );
  sg13g2_a21oi_1 _12380_ (
    .A1(_01445_),
    .A2(_01231_),
    .B1(_02096_),
    .Y(_02098_)
  );
  sg13g2_o21ai_1 _12381_ (
    .A1(_00910_),
    .A2(_02093_),
    .B1(_02098_),
    .Y(_02099_)
  );
  sg13g2_nand2_1 _12382_ (
    .A(_00391_),
    .B(_00368_),
    .Y(_02100_)
  );
  sg13g2_a22oi_1 _12383_ (
    .A1(_01747_),
    .A2(_02100_),
    .B1(_00206_),
    .B2(addr_i_8_),
    .Y(_02101_)
  );
  sg13g2_a22oi_1 _12384_ (
    .A1(_00177_),
    .A2(_00789_),
    .B1(_00933_),
    .B2(addr_i_6_),
    .Y(_02102_)
  );
  sg13g2_nor2_1 _12385_ (
    .A(_03446_),
    .B(_07061_),
    .Y(_02103_)
  );
  sg13g2_nor2_1 _12386_ (
    .A(addr_i_4_),
    .B(_02103_),
    .Y(_02104_)
  );
  sg13g2_buf_1 _12387_ (
    .A(_00535_),
    .X(_02105_)
  );
  sg13g2_o21ai_1 _12388_ (
    .A1(_01194_),
    .A2(_02104_),
    .B1(_02105_),
    .Y(_02106_)
  );
  sg13g2_buf_1 _12389_ (
    .A(_00583_),
    .X(_02107_)
  );
  sg13g2_nand3_1 _12390_ (
    .A(addr_i_2_),
    .B(_04063_),
    .C(_01588_),
    .Y(_02109_)
  );
  sg13g2_a221oi_1 _12391_ (
    .A1(_02107_),
    .A2(_00368_),
    .B1(_02109_),
    .B2(_04981_),
    .C1(_03820_),
    .Y(_02110_)
  );
  sg13g2_a21oi_1 _12392_ (
    .A1(_02102_),
    .A2(_02106_),
    .B1(_02110_),
    .Y(_02111_)
  );
  sg13g2_a221oi_1 _12393_ (
    .A1(addr_i_8_),
    .A2(_02099_),
    .B1(_02101_),
    .B2(_02111_),
    .C1(_00108_),
    .Y(_02112_)
  );
  sg13g2_o21ai_1 _12394_ (
    .A1(_02261_),
    .A2(_01474_),
    .B1(addr_i_6_),
    .Y(_02113_)
  );
  sg13g2_a22oi_1 _12395_ (
    .A1(_01519_),
    .A2(_00770_),
    .B1(_04683_),
    .B2(_00588_),
    .Y(_02114_)
  );
  sg13g2_a21oi_1 _12396_ (
    .A1(addr_i_2_),
    .A2(_05424_),
    .B1(_04086_),
    .Y(_02115_)
  );
  sg13g2_o21ai_1 _12397_ (
    .A1(addr_i_3_),
    .A2(_02115_),
    .B1(_01649_),
    .Y(_02116_)
  );
  sg13g2_a221oi_1 _12398_ (
    .A1(_00861_),
    .A2(_00862_),
    .B1(_02116_),
    .B2(addr_i_4_),
    .C1(_01049_),
    .Y(_02117_)
  );
  sg13g2_nor2_1 _12399_ (
    .A(addr_i_4_),
    .B(_00242_),
    .Y(_02118_)
  );
  sg13g2_o21ai_1 _12400_ (
    .A1(_09226_),
    .A2(_02118_),
    .B1(_00322_),
    .Y(_02120_)
  );
  sg13g2_o21ai_1 _12401_ (
    .A1(_00165_),
    .A2(_03864_),
    .B1(_01537_),
    .Y(_02121_)
  );
  sg13g2_a22oi_1 _12402_ (
    .A1(_00700_),
    .A2(_05280_),
    .B1(_01424_),
    .B2(_02121_),
    .Y(_02122_)
  );
  sg13g2_nor2_1 _12403_ (
    .A(addr_i_3_),
    .B(_03413_),
    .Y(_02123_)
  );
  sg13g2_a21oi_1 _12404_ (
    .A1(_09371_),
    .A2(_01768_),
    .B1(_02086_),
    .Y(_02124_)
  );
  sg13g2_o21ai_1 _12405_ (
    .A1(_02123_),
    .A2(_02124_),
    .B1(addr_i_4_),
    .Y(_02125_)
  );
  sg13g2_nor2_1 _12406_ (
    .A(_00435_),
    .B(_02207_),
    .Y(_02126_)
  );
  sg13g2_o21ai_1 _12407_ (
    .A1(_04782_),
    .A2(_02126_),
    .B1(_05302_),
    .Y(_02127_)
  );
  sg13g2_nand4_1 _12408_ (
    .A(_02120_),
    .B(_02122_),
    .C(_02125_),
    .D(_02127_),
    .Y(_02128_)
  );
  sg13g2_o21ai_1 _12409_ (
    .A1(_08674_),
    .A2(_02117_),
    .B1(_02128_),
    .Y(_02129_)
  );
  sg13g2_a22oi_1 _12410_ (
    .A1(_02113_),
    .A2(_02114_),
    .B1(_02129_),
    .B2(_01452_),
    .Y(_02131_)
  );
  sg13g2_a22oi_1 _12411_ (
    .A1(_00773_),
    .A2(_02087_),
    .B1(_02112_),
    .B2(_02131_),
    .Y(_02132_)
  );
  sg13g2_o21ai_1 _12412_ (
    .A1(_01211_),
    .A2(_02062_),
    .B1(_02132_),
    .Y(_02133_)
  );
  sg13g2_nand2_1 _12413_ (
    .A(addr_i_2_),
    .B(_02283_),
    .Y(_02134_)
  );
  sg13g2_nand2_1 _12414_ (
    .A(_08930_),
    .B(_02134_),
    .Y(_02135_)
  );
  sg13g2_buf_1 _12415_ (
    .A(_00964_),
    .X(_02136_)
  );
  sg13g2_a21oi_1 _12416_ (
    .A1(_06375_),
    .A2(_02136_),
    .B1(_01125_),
    .Y(_02137_)
  );
  sg13g2_a21oi_1 _12417_ (
    .A1(addr_i_4_),
    .A2(_00098_),
    .B1(_02137_),
    .Y(_02138_)
  );
  sg13g2_o21ai_1 _12418_ (
    .A1(addr_i_4_),
    .A2(_02135_),
    .B1(_02138_),
    .Y(_02139_)
  );
  sg13g2_o21ai_1 _12419_ (
    .A1(_01869_),
    .A2(_01966_),
    .B1(addr_i_2_),
    .Y(_02140_)
  );
  sg13g2_a21oi_1 _12420_ (
    .A1(_01594_),
    .A2(_02140_),
    .B1(addr_i_3_),
    .Y(_02142_)
  );
  sg13g2_nor2_1 _12421_ (
    .A(_00030_),
    .B(_01581_),
    .Y(_02143_)
  );
  sg13g2_o21ai_1 _12422_ (
    .A1(_00597_),
    .A2(_02143_),
    .B1(addr_i_7_),
    .Y(_02144_)
  );
  sg13g2_o21ai_1 _12423_ (
    .A1(_01837_),
    .A2(_00257_),
    .B1(addr_i_4_),
    .Y(_02145_)
  );
  sg13g2_nand3_1 _12424_ (
    .A(addr_i_8_),
    .B(_02144_),
    .C(_02145_),
    .Y(_02146_)
  );
  sg13g2_a22oi_1 _12425_ (
    .A1(addr_i_3_),
    .A2(_02139_),
    .B1(_02142_),
    .B2(_02146_),
    .Y(_02147_)
  );
  sg13g2_o21ai_1 _12426_ (
    .A1(addr_i_3_),
    .A2(_01966_),
    .B1(_01152_),
    .Y(_02148_)
  );
  sg13g2_nand2_1 _12427_ (
    .A(_05346_),
    .B(_05225_),
    .Y(_02149_)
  );
  sg13g2_nand2_1 _12428_ (
    .A(_00664_),
    .B(_00635_),
    .Y(_02150_)
  );
  sg13g2_a21oi_1 _12429_ (
    .A1(_02149_),
    .A2(_02150_),
    .B1(_01095_),
    .Y(_02151_)
  );
  sg13g2_nor3_1 _12430_ (
    .A(addr_i_7_),
    .B(addr_i_6_),
    .C(addr_i_5_),
    .Y(_02153_)
  );
  sg13g2_buf_1 _12431_ (
    .A(_02153_),
    .X(_02154_)
  );
  sg13g2_a21oi_1 _12432_ (
    .A1(_00298_),
    .A2(_02154_),
    .B1(_00227_),
    .Y(_02155_)
  );
  sg13g2_nand2_1 _12433_ (
    .A(addr_i_4_),
    .B(_09050_),
    .Y(_02156_)
  );
  sg13g2_a21o_1 _12434_ (
    .A1(_00655_),
    .A2(_02156_),
    .B1(addr_i_2_),
    .X(_02157_)
  );
  sg13g2_o21ai_1 _12435_ (
    .A1(_00047_),
    .A2(_02155_),
    .B1(_02157_),
    .Y(_02158_)
  );
  sg13g2_a22oi_1 _12436_ (
    .A1(_00500_),
    .A2(_02148_),
    .B1(_02151_),
    .B2(_02158_),
    .Y(_02159_)
  );
  sg13g2_o21ai_1 _12437_ (
    .A1(addr_i_8_),
    .A2(_02159_),
    .B1(_09326_),
    .Y(_02160_)
  );
  sg13g2_and2_1 _12438_ (
    .A(_04450_),
    .B(_01765_),
    .X(_02161_)
  );
  sg13g2_a22oi_1 _12439_ (
    .A1(addr_i_3_),
    .A2(_00400_),
    .B1(_00644_),
    .B2(_02161_),
    .Y(_02162_)
  );
  sg13g2_nor2_1 _12440_ (
    .A(addr_i_2_),
    .B(_02162_),
    .Y(_02164_)
  );
  sg13g2_buf_1 _12441_ (
    .A(_01084_),
    .X(_02165_)
  );
  sg13g2_nand2_1 _12442_ (
    .A(_00923_),
    .B(_01352_),
    .Y(_02166_)
  );
  sg13g2_nand2_1 _12443_ (
    .A(_04373_),
    .B(_02166_),
    .Y(_02167_)
  );
  sg13g2_nand2_1 _12444_ (
    .A(_02165_),
    .B(_02167_),
    .Y(_02168_)
  );
  sg13g2_o21ai_1 _12445_ (
    .A1(_02164_),
    .A2(_02168_),
    .B1(addr_i_7_),
    .Y(_02169_)
  );
  sg13g2_nor2_1 _12446_ (
    .A(_00586_),
    .B(_00938_),
    .Y(_02170_)
  );
  sg13g2_nor2_1 _12447_ (
    .A(addr_i_3_),
    .B(_09371_),
    .Y(_02171_)
  );
  sg13g2_nor4_1 _12448_ (
    .A(_01292_),
    .B(_02170_),
    .C(_01863_),
    .D(_02171_),
    .Y(_02172_)
  );
  sg13g2_nand2_1 _12449_ (
    .A(_04418_),
    .B(_00327_),
    .Y(_02173_)
  );
  sg13g2_a21oi_1 _12450_ (
    .A1(_02173_),
    .A2(_00258_),
    .B1(addr_i_7_),
    .Y(_02175_)
  );
  sg13g2_o21ai_1 _12451_ (
    .A1(addr_i_4_),
    .A2(_02172_),
    .B1(_02175_),
    .Y(_02176_)
  );
  sg13g2_nand3_1 _12452_ (
    .A(addr_i_8_),
    .B(_02169_),
    .C(_02176_),
    .Y(_02177_)
  );
  sg13g2_nand2_1 _12453_ (
    .A(addr_i_6_),
    .B(_04650_),
    .Y(_02178_)
  );
  sg13g2_buf_1 _12454_ (
    .A(_02178_),
    .X(_02179_)
  );
  sg13g2_nor2_1 _12455_ (
    .A(_02602_),
    .B(_00238_),
    .Y(_02180_)
  );
  sg13g2_nor2_1 _12456_ (
    .A(addr_i_2_),
    .B(_06209_),
    .Y(_02181_)
  );
  sg13g2_nor2_1 _12457_ (
    .A(addr_i_3_),
    .B(_02181_),
    .Y(_02182_)
  );
  sg13g2_nor3_1 _12458_ (
    .A(_02179_),
    .B(_02180_),
    .C(_02182_),
    .Y(_02183_)
  );
  sg13g2_nor2_1 _12459_ (
    .A(_05424_),
    .B(_03106_),
    .Y(_02184_)
  );
  sg13g2_a21oi_1 _12460_ (
    .A1(_00408_),
    .A2(_01087_),
    .B1(_04041_),
    .Y(_02186_)
  );
  sg13g2_buf_1 _12461_ (
    .A(_00864_),
    .X(_02187_)
  );
  sg13g2_a21oi_1 _12462_ (
    .A1(_00441_),
    .A2(_02187_),
    .B1(addr_i_3_),
    .Y(_02188_)
  );
  sg13g2_nor2_1 _12463_ (
    .A(_02186_),
    .B(_02188_),
    .Y(_02189_)
  );
  sg13g2_o21ai_1 _12464_ (
    .A1(_01169_),
    .A2(_02184_),
    .B1(_02189_),
    .Y(_02190_)
  );
  sg13g2_buf_1 _12465_ (
    .A(_02031_),
    .X(_02191_)
  );
  sg13g2_a22oi_1 _12466_ (
    .A1(addr_i_3_),
    .A2(_02191_),
    .B1(_01184_),
    .B2(_04661_),
    .Y(_02192_)
  );
  sg13g2_nand2b_1 _12467_ (
    .A_N(_02192_),
    .B(addr_i_9_),
    .Y(_02193_)
  );
  sg13g2_a221oi_1 _12468_ (
    .A1(_00845_),
    .A2(_02183_),
    .B1(_02190_),
    .B2(_01633_),
    .C1(_02193_),
    .Y(_02194_)
  );
  sg13g2_a21oi_1 _12469_ (
    .A1(_02177_),
    .A2(_02194_),
    .B1(addr_i_10_),
    .Y(_02195_)
  );
  sg13g2_o21ai_1 _12470_ (
    .A1(_02147_),
    .A2(_02160_),
    .B1(_02195_),
    .Y(_02197_)
  );
  sg13g2_nor3_1 _12471_ (
    .A(addr_i_2_),
    .B(_05169_),
    .C(_01856_),
    .Y(_02198_)
  );
  sg13g2_or2_1 _12472_ (
    .A(_00100_),
    .B(_02198_),
    .X(_02199_)
  );
  sg13g2_nor2_1 _12473_ (
    .A(_08089_),
    .B(_04749_),
    .Y(_02200_)
  );
  sg13g2_o21ai_1 _12474_ (
    .A1(_00104_),
    .A2(_02200_),
    .B1(_00138_),
    .Y(_02201_)
  );
  sg13g2_a22oi_1 _12475_ (
    .A1(addr_i_4_),
    .A2(_02199_),
    .B1(_02201_),
    .B2(_00701_),
    .Y(_02202_)
  );
  sg13g2_buf_1 _12476_ (
    .A(_03632_),
    .X(_02203_)
  );
  sg13g2_a21oi_1 _12477_ (
    .A1(addr_i_5_),
    .A2(_00025_),
    .B1(_00260_),
    .Y(_02204_)
  );
  sg13g2_nor3_1 _12478_ (
    .A(addr_i_3_),
    .B(_02203_),
    .C(_02204_),
    .Y(_02205_)
  );
  sg13g2_nor2_1 _12479_ (
    .A(addr_i_3_),
    .B(_01495_),
    .Y(_02206_)
  );
  sg13g2_o21ai_1 _12480_ (
    .A1(_01739_),
    .A2(_02206_),
    .B1(addr_i_6_),
    .Y(_02208_)
  );
  sg13g2_o21ai_1 _12481_ (
    .A1(_02202_),
    .A2(_02205_),
    .B1(_02208_),
    .Y(_02209_)
  );
  sg13g2_nor3_1 _12482_ (
    .A(addr_i_2_),
    .B(addr_i_7_),
    .C(_08056_),
    .Y(_02210_)
  );
  sg13g2_a21oi_1 _12483_ (
    .A1(_00476_),
    .A2(_01815_),
    .B1(addr_i_3_),
    .Y(_02211_)
  );
  sg13g2_o21ai_1 _12484_ (
    .A1(_02210_),
    .A2(_02211_),
    .B1(addr_i_6_),
    .Y(_02212_)
  );
  sg13g2_buf_1 _12485_ (
    .A(_02558_),
    .X(_02213_)
  );
  sg13g2_nand2_1 _12486_ (
    .A(_02213_),
    .B(_00104_),
    .Y(_02214_)
  );
  sg13g2_nor2_1 _12487_ (
    .A(addr_i_3_),
    .B(_04384_),
    .Y(_02215_)
  );
  sg13g2_a22oi_1 _12488_ (
    .A1(addr_i_2_),
    .A2(_02214_),
    .B1(_02215_),
    .B2(_05645_),
    .Y(_02216_)
  );
  sg13g2_o21ai_1 _12489_ (
    .A1(_01064_),
    .A2(_01138_),
    .B1(addr_i_3_),
    .Y(_02217_)
  );
  sg13g2_nand4_1 _12490_ (
    .A(addr_i_8_),
    .B(_02212_),
    .C(_02216_),
    .D(_02217_),
    .Y(_02219_)
  );
  sg13g2_o21ai_1 _12491_ (
    .A1(addr_i_8_),
    .A2(_02209_),
    .B1(_02219_),
    .Y(_02220_)
  );
  sg13g2_buf_1 _12492_ (
    .A(_00108_),
    .X(_02221_)
  );
  sg13g2_nand2_1 _12493_ (
    .A(_00148_),
    .B(_00873_),
    .Y(_02222_)
  );
  sg13g2_a22oi_1 _12494_ (
    .A1(addr_i_2_),
    .A2(_02222_),
    .B1(_03720_),
    .B2(_07614_),
    .Y(_02223_)
  );
  sg13g2_nor3_1 _12495_ (
    .A(_00726_),
    .B(addr_i_5_),
    .C(_00298_),
    .Y(_02224_)
  );
  sg13g2_o21ai_1 _12496_ (
    .A1(_04683_),
    .A2(_02224_),
    .B1(addr_i_6_),
    .Y(_02225_)
  );
  sg13g2_a21oi_1 _12497_ (
    .A1(addr_i_5_),
    .A2(_05546_),
    .B1(_00347_),
    .Y(_02226_)
  );
  sg13g2_o21ai_1 _12498_ (
    .A1(_00322_),
    .A2(_02226_),
    .B1(addr_i_6_),
    .Y(_02227_)
  );
  sg13g2_a21oi_1 _12499_ (
    .A1(_00736_),
    .A2(_09415_),
    .B1(addr_i_3_),
    .Y(_02228_)
  );
  sg13g2_nor2_1 _12500_ (
    .A(_00550_),
    .B(_01652_),
    .Y(_02230_)
  );
  sg13g2_nor2_1 _12501_ (
    .A(addr_i_4_),
    .B(_02230_),
    .Y(_02231_)
  );
  sg13g2_nor2_1 _12502_ (
    .A(_02228_),
    .B(_02231_),
    .Y(_02232_)
  );
  sg13g2_a21oi_1 _12503_ (
    .A1(_02227_),
    .A2(_02232_),
    .B1(_00802_),
    .Y(_02233_)
  );
  sg13g2_nand2_1 _12504_ (
    .A(_04429_),
    .B(_03314_),
    .Y(_02234_)
  );
  sg13g2_a22oi_1 _12505_ (
    .A1(addr_i_5_),
    .A2(_02234_),
    .B1(_00132_),
    .B2(_00110_),
    .Y(_02235_)
  );
  sg13g2_or2_1 _12506_ (
    .A(_05546_),
    .B(_00299_),
    .X(_02236_)
  );
  sg13g2_o21ai_1 _12507_ (
    .A1(_03281_),
    .A2(_02235_),
    .B1(_02236_),
    .Y(_02237_)
  );
  sg13g2_nor2_1 _12508_ (
    .A(addr_i_2_),
    .B(_02360_),
    .Y(_02238_)
  );
  sg13g2_a21oi_1 _12509_ (
    .A1(_00050_),
    .A2(_00660_),
    .B1(_00065_),
    .Y(_02239_)
  );
  sg13g2_nor2_1 _12510_ (
    .A(_08885_),
    .B(_07746_),
    .Y(_02241_)
  );
  sg13g2_nor2_1 _12511_ (
    .A(_09127_),
    .B(_02241_),
    .Y(_02242_)
  );
  sg13g2_nor4_1 _12512_ (
    .A(addr_i_3_),
    .B(_02238_),
    .C(_02239_),
    .D(_02242_),
    .Y(_02243_)
  );
  sg13g2_o21ai_1 _12513_ (
    .A1(_00695_),
    .A2(_01673_),
    .B1(addr_i_8_),
    .Y(_02244_)
  );
  sg13g2_a221oi_1 _12514_ (
    .A1(addr_i_3_),
    .A2(_02237_),
    .B1(_01967_),
    .B2(_02243_),
    .C1(_02244_),
    .Y(_02245_)
  );
  sg13g2_a22oi_1 _12515_ (
    .A1(_02223_),
    .A2(_02225_),
    .B1(_02233_),
    .B2(_02245_),
    .Y(_02246_)
  );
  sg13g2_nor2_1 _12516_ (
    .A(_02221_),
    .B(_02246_),
    .Y(_02247_)
  );
  sg13g2_a22oi_1 _12517_ (
    .A1(_01176_),
    .A2(_02220_),
    .B1(_02247_),
    .B2(_03040_),
    .Y(_02248_)
  );
  sg13g2_a221oi_1 _12518_ (
    .A1(_01640_),
    .A2(_02133_),
    .B1(_02197_),
    .B2(_02248_),
    .C1(addr_i_12_),
    .Y(_02249_)
  );
  sg13g2_a21o_1 _12519_ (
    .A1(addr_i_12_),
    .A2(_02044_),
    .B1(_02249_),
    .X(data_o_14_)
  );
  sg13g2_buf_1 _12520_ (
    .A(_02996_),
    .X(_02251_)
  );
  sg13g2_o21ai_1 _12521_ (
    .A1(_02744_),
    .A2(_00754_),
    .B1(_02854_),
    .Y(_02252_)
  );
  sg13g2_o21ai_1 _12522_ (
    .A1(_06927_),
    .A2(_00977_),
    .B1(addr_i_3_),
    .Y(_02253_)
  );
  sg13g2_or3_1 _12523_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .C(addr_i_7_),
    .X(_02254_)
  );
  sg13g2_a21oi_1 _12524_ (
    .A1(_03424_),
    .A2(_02254_),
    .B1(_08254_),
    .Y(_02255_)
  );
  sg13g2_nor2_1 _12525_ (
    .A(_04307_),
    .B(_02255_),
    .Y(_02256_)
  );
  sg13g2_buf_1 _12526_ (
    .A(_06375_),
    .X(_02257_)
  );
  sg13g2_a21oi_1 _12527_ (
    .A1(_02253_),
    .A2(_02256_),
    .B1(_02257_),
    .Y(_02258_)
  );
  sg13g2_a21oi_1 _12528_ (
    .A1(addr_i_7_),
    .A2(_02252_),
    .B1(_02258_),
    .Y(_02259_)
  );
  sg13g2_nor2_1 _12529_ (
    .A(_06706_),
    .B(_02259_),
    .Y(_02260_)
  );
  sg13g2_o21ai_1 _12530_ (
    .A1(addr_i_6_),
    .A2(_00415_),
    .B1(addr_i_3_),
    .Y(_02262_)
  );
  sg13g2_o21ai_1 _12531_ (
    .A1(_00159_),
    .A2(_00536_),
    .B1(addr_i_4_),
    .Y(_02263_)
  );
  sg13g2_nor2_1 _12532_ (
    .A(addr_i_4_),
    .B(_00923_),
    .Y(_02264_)
  );
  sg13g2_buf_1 _12533_ (
    .A(_02264_),
    .X(_02265_)
  );
  sg13g2_o21ai_1 _12534_ (
    .A1(_02265_),
    .A2(_01660_),
    .B1(_07149_),
    .Y(_02266_)
  );
  sg13g2_nand3_1 _12535_ (
    .A(_02262_),
    .B(_02263_),
    .C(_02266_),
    .Y(_02267_)
  );
  sg13g2_buf_1 _12536_ (
    .A(_06563_),
    .X(_02268_)
  );
  sg13g2_nor3_1 _12537_ (
    .A(_00046_),
    .B(addr_i_2_),
    .C(_09226_),
    .Y(_02269_)
  );
  sg13g2_o21ai_1 _12538_ (
    .A1(_02268_),
    .A2(_02269_),
    .B1(addr_i_4_),
    .Y(_02270_)
  );
  sg13g2_buf_1 _12539_ (
    .A(_01067_),
    .X(_02271_)
  );
  sg13g2_nand2_1 _12540_ (
    .A(_04650_),
    .B(_01125_),
    .Y(_02273_)
  );
  sg13g2_a21oi_1 _12541_ (
    .A1(_02271_),
    .A2(_00797_),
    .B1(_02273_),
    .Y(_02274_)
  );
  sg13g2_nor2_1 _12542_ (
    .A(_02470_),
    .B(_07724_),
    .Y(_02275_)
  );
  sg13g2_nor3_1 _12543_ (
    .A(_01616_),
    .B(_01285_),
    .C(_02275_),
    .Y(_02276_)
  );
  sg13g2_buf_1 _12544_ (
    .A(_00744_),
    .X(_02277_)
  );
  sg13g2_nand2_1 _12545_ (
    .A(_06364_),
    .B(_04318_),
    .Y(_02278_)
  );
  sg13g2_a21oi_1 _12546_ (
    .A1(_02277_),
    .A2(_02278_),
    .B1(_00133_),
    .Y(_02279_)
  );
  sg13g2_a221oi_1 _12547_ (
    .A1(_02270_),
    .A2(_02274_),
    .B1(_02276_),
    .B2(_02279_),
    .C1(addr_i_9_),
    .Y(_02280_)
  );
  sg13g2_o21ai_1 _12548_ (
    .A1(_01082_),
    .A2(_02267_),
    .B1(_02280_),
    .Y(_02281_)
  );
  sg13g2_o21ai_1 _12549_ (
    .A1(_01112_),
    .A2(_09183_),
    .B1(_01528_),
    .Y(_02282_)
  );
  sg13g2_o21ai_1 _12550_ (
    .A1(_00534_),
    .A2(_00559_),
    .B1(addr_i_3_),
    .Y(_02284_)
  );
  sg13g2_o21ai_1 _12551_ (
    .A1(_08896_),
    .A2(_09348_),
    .B1(addr_i_4_),
    .Y(_02285_)
  );
  sg13g2_nand4_1 _12552_ (
    .A(_01354_),
    .B(_02282_),
    .C(_02284_),
    .D(_02285_),
    .Y(_02286_)
  );
  sg13g2_buf_1 _12553_ (
    .A(_00260_),
    .X(_02287_)
  );
  sg13g2_o21ai_1 _12554_ (
    .A1(addr_i_4_),
    .A2(_00990_),
    .B1(_02287_),
    .Y(_02288_)
  );
  sg13g2_nor2_1 _12555_ (
    .A(addr_i_6_),
    .B(_05943_),
    .Y(_02289_)
  );
  sg13g2_nand2_1 _12556_ (
    .A(_06054_),
    .B(_01697_),
    .Y(_02290_)
  );
  sg13g2_o21ai_1 _12557_ (
    .A1(addr_i_5_),
    .A2(_02289_),
    .B1(_02290_),
    .Y(_02291_)
  );
  sg13g2_a22oi_1 _12558_ (
    .A1(addr_i_3_),
    .A2(_02288_),
    .B1(_02291_),
    .B2(addr_i_7_),
    .Y(_02292_)
  );
  sg13g2_nand3_1 _12559_ (
    .A(_00080_),
    .B(_09499_),
    .C(_01749_),
    .Y(_02293_)
  );
  sg13g2_nand2_1 _12560_ (
    .A(_00113_),
    .B(_02293_),
    .Y(_02295_)
  );
  sg13g2_a22oi_1 _12561_ (
    .A1(addr_i_7_),
    .A2(_02286_),
    .B1(_02292_),
    .B2(_02295_),
    .Y(_02296_)
  );
  sg13g2_buf_1 _12562_ (
    .A(_05546_),
    .X(_02297_)
  );
  sg13g2_xnor2_1 _12563_ (
    .A(_06154_),
    .B(_05535_),
    .Y(_02298_)
  );
  sg13g2_nand2_1 _12564_ (
    .A(_02297_),
    .B(_02298_),
    .Y(_02299_)
  );
  sg13g2_nand3_1 _12565_ (
    .A(addr_i_3_),
    .B(_00651_),
    .C(_00173_),
    .Y(_02300_)
  );
  sg13g2_nand3_1 _12566_ (
    .A(_00485_),
    .B(_00080_),
    .C(_00704_),
    .Y(_02301_)
  );
  sg13g2_a21oi_1 _12567_ (
    .A1(_02300_),
    .A2(_02301_),
    .B1(_00053_),
    .Y(_02302_)
  );
  sg13g2_o21ai_1 _12568_ (
    .A1(_02026_),
    .A2(_00156_),
    .B1(_05247_),
    .Y(_02303_)
  );
  sg13g2_nand2_1 _12569_ (
    .A(addr_i_5_),
    .B(_06840_),
    .Y(_02304_)
  );
  sg13g2_nand3_1 _12570_ (
    .A(_01878_),
    .B(_00314_),
    .C(_02304_),
    .Y(_02306_)
  );
  sg13g2_nand3_1 _12571_ (
    .A(addr_i_8_),
    .B(_02303_),
    .C(_02306_),
    .Y(_02307_)
  );
  sg13g2_a22oi_1 _12572_ (
    .A1(_01892_),
    .A2(_02299_),
    .B1(_02302_),
    .B2(_02307_),
    .Y(_02308_)
  );
  sg13g2_o21ai_1 _12573_ (
    .A1(_02296_),
    .A2(_02308_),
    .B1(addr_i_9_),
    .Y(_02309_)
  );
  sg13g2_o21ai_1 _12574_ (
    .A1(_02260_),
    .A2(_02281_),
    .B1(_02309_),
    .Y(_02310_)
  );
  sg13g2_nand2_1 _12575_ (
    .A(addr_i_10_),
    .B(_02310_),
    .Y(_02311_)
  );
  sg13g2_nand2_1 _12576_ (
    .A(addr_i_6_),
    .B(_00679_),
    .Y(_02312_)
  );
  sg13g2_nand2_1 _12577_ (
    .A(_00343_),
    .B(_02312_),
    .Y(_02313_)
  );
  sg13g2_a21oi_1 _12578_ (
    .A1(_07094_),
    .A2(_02313_),
    .B1(_02271_),
    .Y(_02314_)
  );
  sg13g2_nand2_1 _12579_ (
    .A(_01585_),
    .B(_09494_),
    .Y(_02315_)
  );
  sg13g2_a21oi_1 _12580_ (
    .A1(_01499_),
    .A2(_02315_),
    .B1(addr_i_3_),
    .Y(_02317_)
  );
  sg13g2_o21ai_1 _12581_ (
    .A1(_02314_),
    .A2(_02317_),
    .B1(addr_i_2_),
    .Y(_02318_)
  );
  sg13g2_nand2_1 _12582_ (
    .A(_07105_),
    .B(_03665_),
    .Y(_02319_)
  );
  sg13g2_o21ai_1 _12583_ (
    .A1(addr_i_3_),
    .A2(_09504_),
    .B1(_02319_),
    .Y(_02320_)
  );
  sg13g2_a21oi_1 _12584_ (
    .A1(addr_i_4_),
    .A2(_00678_),
    .B1(_05700_),
    .Y(_02321_)
  );
  sg13g2_nor2_1 _12585_ (
    .A(addr_i_4_),
    .B(_00678_),
    .Y(_02322_)
  );
  sg13g2_nor3_1 _12586_ (
    .A(_01232_),
    .B(_02321_),
    .C(_02322_),
    .Y(_02323_)
  );
  sg13g2_a21oi_1 _12587_ (
    .A1(_04041_),
    .A2(_08254_),
    .B1(_00343_),
    .Y(_02324_)
  );
  sg13g2_nor2_1 _12588_ (
    .A(addr_i_2_),
    .B(_02324_),
    .Y(_02325_)
  );
  sg13g2_a221oi_1 _12589_ (
    .A1(addr_i_5_),
    .A2(_02320_),
    .B1(_02323_),
    .B2(_02325_),
    .C1(addr_i_9_),
    .Y(_02326_)
  );
  sg13g2_a21oi_1 _12590_ (
    .A1(_00343_),
    .A2(_00473_),
    .B1(_07647_),
    .Y(_02328_)
  );
  sg13g2_nor2_1 _12591_ (
    .A(addr_i_5_),
    .B(_05379_),
    .Y(_02329_)
  );
  sg13g2_nor2_1 _12592_ (
    .A(_05281_),
    .B(_01066_),
    .Y(_02330_)
  );
  sg13g2_a22oi_1 _12593_ (
    .A1(addr_i_4_),
    .A2(_02329_),
    .B1(_02330_),
    .B2(_00119_),
    .Y(_02331_)
  );
  sg13g2_o21ai_1 _12594_ (
    .A1(addr_i_3_),
    .A2(_02328_),
    .B1(_02331_),
    .Y(_02332_)
  );
  sg13g2_nor2_1 _12595_ (
    .A(_08166_),
    .B(_03864_),
    .Y(_02333_)
  );
  sg13g2_o21ai_1 _12596_ (
    .A1(_00731_),
    .A2(_01222_),
    .B1(addr_i_9_),
    .Y(_02334_)
  );
  sg13g2_a21o_1 _12597_ (
    .A1(_00150_),
    .A2(_02333_),
    .B1(_02334_),
    .X(_02335_)
  );
  sg13g2_a21oi_1 _12598_ (
    .A1(_09473_),
    .A2(_00783_),
    .B1(_00743_),
    .Y(_02336_)
  );
  sg13g2_o21ai_1 _12599_ (
    .A1(_00100_),
    .A2(_08299_),
    .B1(_00822_),
    .Y(_02337_)
  );
  sg13g2_a21oi_1 _12600_ (
    .A1(_02336_),
    .A2(_02337_),
    .B1(addr_i_4_),
    .Y(_02339_)
  );
  sg13g2_a22oi_1 _12601_ (
    .A1(addr_i_7_),
    .A2(_02332_),
    .B1(_02335_),
    .B2(_02339_),
    .Y(_02340_)
  );
  sg13g2_a22oi_1 _12602_ (
    .A1(_02318_),
    .A2(_02326_),
    .B1(_06706_),
    .B2(_02340_),
    .Y(_02341_)
  );
  sg13g2_nor2_1 _12603_ (
    .A(_00199_),
    .B(_00303_),
    .Y(_02342_)
  );
  sg13g2_buf_1 _12604_ (
    .A(_00064_),
    .X(_02343_)
  );
  sg13g2_buf_1 _12605_ (
    .A(_02343_),
    .X(_02344_)
  );
  sg13g2_nor3_1 _12606_ (
    .A(_02344_),
    .B(_00949_),
    .C(_05600_),
    .Y(_02345_)
  );
  sg13g2_a221oi_1 _12607_ (
    .A1(addr_i_4_),
    .A2(_00317_),
    .B1(_01216_),
    .B2(_00074_),
    .C1(_02345_),
    .Y(_02346_)
  );
  sg13g2_a21oi_1 _12608_ (
    .A1(addr_i_7_),
    .A2(_06873_),
    .B1(_01031_),
    .Y(_02347_)
  );
  sg13g2_nor4_1 _12609_ (
    .A(_00374_),
    .B(addr_i_8_),
    .C(_00087_),
    .D(_02069_),
    .Y(_02348_)
  );
  sg13g2_o21ai_1 _12610_ (
    .A1(_08266_),
    .A2(_02347_),
    .B1(_02348_),
    .Y(_02350_)
  );
  sg13g2_a221oi_1 _12611_ (
    .A1(_01336_),
    .A2(_02342_),
    .B1(_02346_),
    .B2(addr_i_3_),
    .C1(_02350_),
    .Y(_02351_)
  );
  sg13g2_a21oi_1 _12612_ (
    .A1(addr_i_5_),
    .A2(_00194_),
    .B1(_01159_),
    .Y(_02352_)
  );
  sg13g2_o21ai_1 _12613_ (
    .A1(addr_i_3_),
    .A2(_02352_),
    .B1(_00317_),
    .Y(_02353_)
  );
  sg13g2_nand2_1 _12614_ (
    .A(addr_i_2_),
    .B(_02353_),
    .Y(_02354_)
  );
  sg13g2_a21oi_1 _12615_ (
    .A1(_00185_),
    .A2(_09508_),
    .B1(addr_i_2_),
    .Y(_02355_)
  );
  sg13g2_o21ai_1 _12616_ (
    .A1(_00898_),
    .A2(_02355_),
    .B1(_01794_),
    .Y(_02356_)
  );
  sg13g2_o21ai_1 _12617_ (
    .A1(_06950_),
    .A2(_05258_),
    .B1(_00091_),
    .Y(_02357_)
  );
  sg13g2_o21ai_1 _12618_ (
    .A1(_06398_),
    .A2(_00977_),
    .B1(addr_i_4_),
    .Y(_02358_)
  );
  sg13g2_nand2_1 _12619_ (
    .A(_02357_),
    .B(_02358_),
    .Y(_02359_)
  );
  sg13g2_nor2_1 _12620_ (
    .A(_00586_),
    .B(_06077_),
    .Y(_02361_)
  );
  sg13g2_a22oi_1 _12621_ (
    .A1(addr_i_3_),
    .A2(_02359_),
    .B1(_02361_),
    .B2(_00214_),
    .Y(_02362_)
  );
  sg13g2_and3_1 _12622_ (
    .A(_02354_),
    .B(_02356_),
    .C(_02362_),
    .X(_02363_)
  );
  sg13g2_or4_1 _12623_ (
    .A(addr_i_10_),
    .B(_02341_),
    .C(_02351_),
    .D(_02363_),
    .X(_02364_)
  );
  sg13g2_nand3_1 _12624_ (
    .A(_02251_),
    .B(_02311_),
    .C(_02364_),
    .Y(_02365_)
  );
  sg13g2_nor2_1 _12625_ (
    .A(_00191_),
    .B(_00959_),
    .Y(_02366_)
  );
  sg13g2_a21oi_1 _12626_ (
    .A1(addr_i_7_),
    .A2(_09105_),
    .B1(_02366_),
    .Y(_02367_)
  );
  sg13g2_buf_1 _12627_ (
    .A(_00214_),
    .X(_02368_)
  );
  sg13g2_nor2b_1 _12628_ (
    .A(addr_i_7_),
    .B_N(addr_i_3_),
    .Y(_02369_)
  );
  sg13g2_a22oi_1 _12629_ (
    .A1(_09094_),
    .A2(_00645_),
    .B1(_02369_),
    .B2(_00172_),
    .Y(_02370_)
  );
  sg13g2_nor2_1 _12630_ (
    .A(_02368_),
    .B(_02370_),
    .Y(_02372_)
  );
  sg13g2_o21ai_1 _12631_ (
    .A1(addr_i_6_),
    .A2(_02367_),
    .B1(_02372_),
    .Y(_02373_)
  );
  sg13g2_nor2_1 _12632_ (
    .A(_01160_),
    .B(_00516_),
    .Y(_02374_)
  );
  sg13g2_nor2_1 _12633_ (
    .A(addr_i_7_),
    .B(_02374_),
    .Y(_02375_)
  );
  sg13g2_nor2_1 _12634_ (
    .A(addr_i_3_),
    .B(_09493_),
    .Y(_02376_)
  );
  sg13g2_nor2_1 _12635_ (
    .A(_00401_),
    .B(_00531_),
    .Y(_02377_)
  );
  sg13g2_o21ai_1 _12636_ (
    .A1(_02376_),
    .A2(_02377_),
    .B1(_00123_),
    .Y(_02378_)
  );
  sg13g2_a21oi_1 _12637_ (
    .A1(_02375_),
    .A2(_02378_),
    .B1(_02368_),
    .Y(_02379_)
  );
  sg13g2_nor2_1 _12638_ (
    .A(addr_i_3_),
    .B(_07956_),
    .Y(_02380_)
  );
  sg13g2_o21ai_1 _12639_ (
    .A1(_04683_),
    .A2(_02380_),
    .B1(addr_i_6_),
    .Y(_02381_)
  );
  sg13g2_nand2_1 _12640_ (
    .A(_03446_),
    .B(_05910_),
    .Y(_02383_)
  );
  sg13g2_nor2_1 _12641_ (
    .A(_00047_),
    .B(_02383_),
    .Y(_02384_)
  );
  sg13g2_o21ai_1 _12642_ (
    .A1(_00523_),
    .A2(_02384_),
    .B1(_00068_),
    .Y(_02385_)
  );
  sg13g2_nand3_1 _12643_ (
    .A(addr_i_7_),
    .B(_02381_),
    .C(_02385_),
    .Y(_02386_)
  );
  sg13g2_buf_1 _12644_ (
    .A(_05324_),
    .X(_02387_)
  );
  sg13g2_nor2_1 _12645_ (
    .A(_06530_),
    .B(_03632_),
    .Y(_02388_)
  );
  sg13g2_nor2_1 _12646_ (
    .A(_02387_),
    .B(_02388_),
    .Y(_02389_)
  );
  sg13g2_o21ai_1 _12647_ (
    .A1(_00119_),
    .A2(_02389_),
    .B1(_00068_),
    .Y(_02390_)
  );
  sg13g2_nor2_1 _12648_ (
    .A(_05745_),
    .B(_00516_),
    .Y(_02391_)
  );
  sg13g2_a22oi_1 _12649_ (
    .A1(addr_i_2_),
    .A2(_00905_),
    .B1(_02391_),
    .B2(addr_i_7_),
    .Y(_02392_)
  );
  sg13g2_a22oi_1 _12650_ (
    .A1(_02390_),
    .A2(_02392_),
    .B1(_00386_),
    .B2(_01612_),
    .Y(_02394_)
  );
  sg13g2_nor2_1 _12651_ (
    .A(_05379_),
    .B(_00605_),
    .Y(_02395_)
  );
  sg13g2_a21oi_1 _12652_ (
    .A1(_00780_),
    .A2(_01274_),
    .B1(addr_i_4_),
    .Y(_02396_)
  );
  sg13g2_a21oi_1 _12653_ (
    .A1(addr_i_4_),
    .A2(_00429_),
    .B1(_02396_),
    .Y(_02397_)
  );
  sg13g2_o21ai_1 _12654_ (
    .A1(_07514_),
    .A2(_02395_),
    .B1(_02397_),
    .Y(_02398_)
  );
  sg13g2_a21o_1 _12655_ (
    .A1(addr_i_9_),
    .A2(_02398_),
    .B1(addr_i_10_),
    .X(_02399_)
  );
  sg13g2_a22oi_1 _12656_ (
    .A1(_02379_),
    .A2(_02386_),
    .B1(_02394_),
    .B2(_02399_),
    .Y(_02400_)
  );
  sg13g2_a22oi_1 _12657_ (
    .A1(addr_i_10_),
    .A2(_02373_),
    .B1(_02400_),
    .B2(_00812_),
    .Y(_02401_)
  );
  sg13g2_nor2_1 _12658_ (
    .A(_03051_),
    .B(_02401_),
    .Y(_02402_)
  );
  sg13g2_o21ai_1 _12659_ (
    .A1(addr_i_6_),
    .A2(addr_i_5_),
    .B1(addr_i_7_),
    .Y(_02403_)
  );
  sg13g2_buf_1 _12660_ (
    .A(_02403_),
    .X(_02405_)
  );
  sg13g2_nand2_1 _12661_ (
    .A(_05966_),
    .B(_04926_),
    .Y(_02406_)
  );
  sg13g2_o21ai_1 _12662_ (
    .A1(addr_i_2_),
    .A2(_02405_),
    .B1(_02406_),
    .Y(_02407_)
  );
  sg13g2_a21oi_1 _12663_ (
    .A1(_01221_),
    .A2(_01601_),
    .B1(addr_i_4_),
    .Y(_02408_)
  );
  sg13g2_a22oi_1 _12664_ (
    .A1(addr_i_4_),
    .A2(_02407_),
    .B1(_02408_),
    .B2(_07425_),
    .Y(_02409_)
  );
  sg13g2_nand2_1 _12665_ (
    .A(_02250_),
    .B(_01084_),
    .Y(_02410_)
  );
  sg13g2_nand2_1 _12666_ (
    .A(_08597_),
    .B(_04528_),
    .Y(_02411_)
  );
  sg13g2_o21ai_1 _12667_ (
    .A1(addr_i_7_),
    .A2(_00219_),
    .B1(_02411_),
    .Y(_02412_)
  );
  sg13g2_nand3_1 _12668_ (
    .A(addr_i_7_),
    .B(_02031_),
    .C(_01084_),
    .Y(_02413_)
  );
  sg13g2_a21oi_1 _12669_ (
    .A1(_09475_),
    .A2(_02413_),
    .B1(addr_i_6_),
    .Y(_02414_)
  );
  sg13g2_a22oi_1 _12670_ (
    .A1(addr_i_6_),
    .A2(_02410_),
    .B1(_02412_),
    .B2(_02414_),
    .Y(_02416_)
  );
  sg13g2_mux2_1 _12671_ (
    .A0(_02409_),
    .A1(_02416_),
    .S(_08752_),
    .X(_02417_)
  );
  sg13g2_nor2_1 _12672_ (
    .A(_00384_),
    .B(_00234_),
    .Y(_02418_)
  );
  sg13g2_nor2_1 _12673_ (
    .A(_05722_),
    .B(_02031_),
    .Y(_02419_)
  );
  sg13g2_nor2_1 _12674_ (
    .A(_02371_),
    .B(_00406_),
    .Y(_02420_)
  );
  sg13g2_o21ai_1 _12675_ (
    .A1(_02419_),
    .A2(_02420_),
    .B1(addr_i_3_),
    .Y(_02421_)
  );
  sg13g2_o21ai_1 _12676_ (
    .A1(_02755_),
    .A2(_02418_),
    .B1(_02421_),
    .Y(_02422_)
  );
  sg13g2_nor3_1 _12677_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .C(addr_i_5_),
    .Y(_02423_)
  );
  sg13g2_buf_1 _12678_ (
    .A(_02423_),
    .X(_02424_)
  );
  sg13g2_nor2_1 _12679_ (
    .A(_07757_),
    .B(_02424_),
    .Y(_02425_)
  );
  sg13g2_nand2_1 _12680_ (
    .A(addr_i_7_),
    .B(_00616_),
    .Y(_02427_)
  );
  sg13g2_nor2_1 _12681_ (
    .A(_00030_),
    .B(_07160_),
    .Y(_02428_)
  );
  sg13g2_a21oi_1 _12682_ (
    .A1(_00965_),
    .A2(_02887_),
    .B1(_08741_),
    .Y(_02429_)
  );
  sg13g2_o21ai_1 _12683_ (
    .A1(_02428_),
    .A2(_02429_),
    .B1(addr_i_2_),
    .Y(_02430_)
  );
  sg13g2_o21ai_1 _12684_ (
    .A1(_02425_),
    .A2(_02427_),
    .B1(_02430_),
    .Y(_02431_)
  );
  sg13g2_a22oi_1 _12685_ (
    .A1(_04052_),
    .A2(_02422_),
    .B1(_02431_),
    .B2(addr_i_8_),
    .Y(_02432_)
  );
  sg13g2_a21oi_1 _12686_ (
    .A1(addr_i_8_),
    .A2(_02417_),
    .B1(_02432_),
    .Y(_02433_)
  );
  sg13g2_nand2_1 _12687_ (
    .A(_07967_),
    .B(_00665_),
    .Y(_02434_)
  );
  sg13g2_nand2_1 _12688_ (
    .A(_02191_),
    .B(_08553_),
    .Y(_02435_)
  );
  sg13g2_a21oi_1 _12689_ (
    .A1(_02434_),
    .A2(_02435_),
    .B1(addr_i_3_),
    .Y(_02436_)
  );
  sg13g2_nand2_1 _12690_ (
    .A(addr_i_3_),
    .B(_07724_),
    .Y(_02438_)
  );
  sg13g2_o21ai_1 _12691_ (
    .A1(_00558_),
    .A2(_02438_),
    .B1(_01633_),
    .Y(_02439_)
  );
  sg13g2_nand3_1 _12692_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .C(_06485_),
    .Y(_02440_)
  );
  sg13g2_nor2_1 _12693_ (
    .A(addr_i_4_),
    .B(_07469_),
    .Y(_02441_)
  );
  sg13g2_o21ai_1 _12694_ (
    .A1(_02441_),
    .A2(_01306_),
    .B1(_00347_),
    .Y(_02442_)
  );
  sg13g2_nor2_1 _12695_ (
    .A(addr_i_4_),
    .B(_01965_),
    .Y(_02443_)
  );
  sg13g2_o21ai_1 _12696_ (
    .A1(_01401_),
    .A2(_02443_),
    .B1(addr_i_3_),
    .Y(_02444_)
  );
  sg13g2_nand3_1 _12697_ (
    .A(_02440_),
    .B(_02442_),
    .C(_02444_),
    .Y(_02445_)
  );
  sg13g2_o21ai_1 _12698_ (
    .A1(_02503_),
    .A2(_01735_),
    .B1(addr_i_6_),
    .Y(_02446_)
  );
  sg13g2_a21oi_1 _12699_ (
    .A1(_05689_),
    .A2(_01028_),
    .B1(_08741_),
    .Y(_02447_)
  );
  sg13g2_a21oi_1 _12700_ (
    .A1(addr_i_2_),
    .A2(_03117_),
    .B1(_02447_),
    .Y(_02449_)
  );
  sg13g2_a21oi_1 _12701_ (
    .A1(_02446_),
    .A2(_02449_),
    .B1(_00791_),
    .Y(_02450_)
  );
  sg13g2_nand3_1 _12702_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .C(_04418_),
    .Y(_02451_)
  );
  sg13g2_a21oi_1 _12703_ (
    .A1(_00413_),
    .A2(_02451_),
    .B1(_05711_),
    .Y(_02452_)
  );
  sg13g2_and2_1 _12704_ (
    .A(_00463_),
    .B(_07480_),
    .X(_02453_)
  );
  sg13g2_a21oi_1 _12705_ (
    .A1(addr_i_2_),
    .A2(_07779_),
    .B1(addr_i_4_),
    .Y(_02454_)
  );
  sg13g2_nor4_1 _12706_ (
    .A(_01494_),
    .B(_02452_),
    .C(_02453_),
    .D(_02454_),
    .Y(_02455_)
  );
  sg13g2_a22oi_1 _12707_ (
    .A1(_01666_),
    .A2(_02445_),
    .B1(_02450_),
    .B2(_02455_),
    .Y(_02456_)
  );
  sg13g2_o21ai_1 _12708_ (
    .A1(_02436_),
    .A2(_02439_),
    .B1(_02456_),
    .Y(_02457_)
  );
  sg13g2_mux2_1 _12709_ (
    .A0(_02433_),
    .A1(_02457_),
    .S(_04705_),
    .X(_02458_)
  );
  sg13g2_nor3_1 _12710_ (
    .A(_08156_),
    .B(_00165_),
    .C(_00242_),
    .Y(_02460_)
  );
  sg13g2_o21ai_1 _12711_ (
    .A1(_00897_),
    .A2(_02460_),
    .B1(addr_i_2_),
    .Y(_02461_)
  );
  sg13g2_buf_1 _12712_ (
    .A(_00998_),
    .X(_02462_)
  );
  sg13g2_o21ai_1 _12713_ (
    .A1(_00269_),
    .A2(_01587_),
    .B1(_02462_),
    .Y(_02463_)
  );
  sg13g2_nand3_1 _12714_ (
    .A(_00476_),
    .B(_02461_),
    .C(_02463_),
    .Y(_02464_)
  );
  sg13g2_o21ai_1 _12715_ (
    .A1(_08100_),
    .A2(_00100_),
    .B1(_00719_),
    .Y(_02465_)
  );
  sg13g2_a21oi_1 _12716_ (
    .A1(_08707_),
    .A2(_02465_),
    .B1(addr_i_4_),
    .Y(_02466_)
  );
  sg13g2_buf_1 _12717_ (
    .A(_00671_),
    .X(_02467_)
  );
  sg13g2_a21oi_1 _12718_ (
    .A1(_00476_),
    .A2(_02467_),
    .B1(_00820_),
    .Y(_02468_)
  );
  sg13g2_a22oi_1 _12719_ (
    .A1(addr_i_4_),
    .A2(_02464_),
    .B1(_02466_),
    .B2(_02468_),
    .Y(_02469_)
  );
  sg13g2_buf_1 _12720_ (
    .A(_02360_),
    .X(_02471_)
  );
  sg13g2_buf_1 _12721_ (
    .A(_08564_),
    .X(_02472_)
  );
  sg13g2_nor2_1 _12722_ (
    .A(_02471_),
    .B(_02472_),
    .Y(_02473_)
  );
  sg13g2_nand4_1 _12723_ (
    .A(addr_i_4_),
    .B(_03809_),
    .C(_01581_),
    .D(_01273_),
    .Y(_02474_)
  );
  sg13g2_o21ai_1 _12724_ (
    .A1(_02136_),
    .A2(_00911_),
    .B1(_02474_),
    .Y(_02475_)
  );
  sg13g2_o21ai_1 _12725_ (
    .A1(_02473_),
    .A2(_02475_),
    .B1(addr_i_3_),
    .Y(_02476_)
  );
  sg13g2_o21ai_1 _12726_ (
    .A1(_00484_),
    .A2(_00624_),
    .B1(_00956_),
    .Y(_02477_)
  );
  sg13g2_a21oi_1 _12727_ (
    .A1(_00505_),
    .A2(_02477_),
    .B1(addr_i_3_),
    .Y(_02478_)
  );
  sg13g2_buf_1 _12728_ (
    .A(_01625_),
    .X(_02479_)
  );
  sg13g2_a21oi_1 _12729_ (
    .A1(_00582_),
    .A2(_02479_),
    .B1(addr_i_6_),
    .Y(_02480_)
  );
  sg13g2_nor2_1 _12730_ (
    .A(_02478_),
    .B(_02480_),
    .Y(_02482_)
  );
  sg13g2_a21oi_1 _12731_ (
    .A1(_02476_),
    .A2(_02482_),
    .B1(addr_i_8_),
    .Y(_02483_)
  );
  sg13g2_a21oi_1 _12732_ (
    .A1(addr_i_8_),
    .A2(_02469_),
    .B1(_02483_),
    .Y(_02484_)
  );
  sg13g2_o21ai_1 _12733_ (
    .A1(_05025_),
    .A2(_07879_),
    .B1(_04119_),
    .Y(_02485_)
  );
  sg13g2_nor2_1 _12734_ (
    .A(_05324_),
    .B(_09493_),
    .Y(_02486_)
  );
  sg13g2_o21ai_1 _12735_ (
    .A1(_00234_),
    .A2(_02486_),
    .B1(addr_i_2_),
    .Y(_02487_)
  );
  sg13g2_nand3_1 _12736_ (
    .A(_01203_),
    .B(_02485_),
    .C(_02487_),
    .Y(_02488_)
  );
  sg13g2_o21ai_1 _12737_ (
    .A1(_08896_),
    .A2(_01276_),
    .B1(addr_i_4_),
    .Y(_02489_)
  );
  sg13g2_nor2_1 _12738_ (
    .A(addr_i_3_),
    .B(_07746_),
    .Y(_02490_)
  );
  sg13g2_a221oi_1 _12739_ (
    .A1(_08177_),
    .A2(_02489_),
    .B1(_02490_),
    .B2(_01050_),
    .C1(_00778_),
    .Y(_02491_)
  );
  sg13g2_a21o_1 _12740_ (
    .A1(_04052_),
    .A2(_02488_),
    .B1(_02491_),
    .X(_02493_)
  );
  sg13g2_nand2_1 _12741_ (
    .A(_02343_),
    .B(_00498_),
    .Y(_02494_)
  );
  sg13g2_nand3_1 _12742_ (
    .A(_00022_),
    .B(_00429_),
    .C(_02494_),
    .Y(_02495_)
  );
  sg13g2_nand2_1 _12743_ (
    .A(addr_i_3_),
    .B(_04075_),
    .Y(_02496_)
  );
  sg13g2_nand2_1 _12744_ (
    .A(_00354_),
    .B(_01179_),
    .Y(_02497_)
  );
  sg13g2_nor2_1 _12745_ (
    .A(_06386_),
    .B(_01000_),
    .Y(_02498_)
  );
  sg13g2_nand3_1 _12746_ (
    .A(_02496_),
    .B(_02497_),
    .C(_02498_),
    .Y(_02499_)
  );
  sg13g2_nor2_1 _12747_ (
    .A(addr_i_3_),
    .B(_02241_),
    .Y(_02500_)
  );
  sg13g2_nor2_1 _12748_ (
    .A(addr_i_6_),
    .B(_01011_),
    .Y(_02501_)
  );
  sg13g2_o21ai_1 _12749_ (
    .A1(_01187_),
    .A2(_02500_),
    .B1(_02501_),
    .Y(_02502_)
  );
  sg13g2_nand4_1 _12750_ (
    .A(addr_i_9_),
    .B(_02495_),
    .C(_02499_),
    .D(_02502_),
    .Y(_02504_)
  );
  sg13g2_nand2_1 _12751_ (
    .A(addr_i_6_),
    .B(_00079_),
    .Y(_02505_)
  );
  sg13g2_a21oi_1 _12752_ (
    .A1(_09483_),
    .A2(_02505_),
    .B1(_02271_),
    .Y(_02506_)
  );
  sg13g2_nand2_1 _12753_ (
    .A(_00736_),
    .B(_03139_),
    .Y(_02507_)
  );
  sg13g2_a21oi_1 _12754_ (
    .A1(_01367_),
    .A2(_02507_),
    .B1(addr_i_3_),
    .Y(_02508_)
  );
  sg13g2_nor4_1 _12755_ (
    .A(_07403_),
    .B(_01380_),
    .C(_02506_),
    .D(_02508_),
    .Y(_02509_)
  );
  sg13g2_a22oi_1 _12756_ (
    .A1(_01151_),
    .A2(_02493_),
    .B1(_02504_),
    .B2(_02509_),
    .Y(_02510_)
  );
  sg13g2_a22oi_1 _12757_ (
    .A1(_09326_),
    .A2(_02484_),
    .B1(_02510_),
    .B2(addr_i_12_),
    .Y(_02511_)
  );
  sg13g2_a21o_1 _12758_ (
    .A1(addr_i_12_),
    .A2(_02458_),
    .B1(_02511_),
    .X(_02512_)
  );
  sg13g2_buf_1 _12759_ (
    .A(_08520_),
    .X(_02513_)
  );
  sg13g2_nand2_1 _12760_ (
    .A(_00930_),
    .B(_02513_),
    .Y(_02515_)
  );
  sg13g2_a22oi_1 _12761_ (
    .A1(addr_i_5_),
    .A2(_02515_),
    .B1(_02203_),
    .B2(addr_i_2_),
    .Y(_02516_)
  );
  sg13g2_nand2_1 _12762_ (
    .A(addr_i_2_),
    .B(_00316_),
    .Y(_02517_)
  );
  sg13g2_a21oi_1 _12763_ (
    .A1(_00070_),
    .A2(_00695_),
    .B1(addr_i_5_),
    .Y(_02518_)
  );
  sg13g2_nor2_1 _12764_ (
    .A(_02517_),
    .B(_02518_),
    .Y(_02519_)
  );
  sg13g2_o21ai_1 _12765_ (
    .A1(_02516_),
    .A2(_02519_),
    .B1(addr_i_3_),
    .Y(_02520_)
  );
  sg13g2_nand3_1 _12766_ (
    .A(addr_i_5_),
    .B(_00492_),
    .C(_00414_),
    .Y(_02521_)
  );
  sg13g2_nand2_1 _12767_ (
    .A(_08232_),
    .B(_02521_),
    .Y(_02522_)
  );
  sg13g2_nor3_1 _12768_ (
    .A(addr_i_5_),
    .B(_06927_),
    .C(_09473_),
    .Y(_02523_)
  );
  sg13g2_a22oi_1 _12769_ (
    .A1(addr_i_5_),
    .A2(_09492_),
    .B1(_02523_),
    .B2(addr_i_2_),
    .Y(_02524_)
  );
  sg13g2_a22oi_1 _12770_ (
    .A1(_00084_),
    .A2(_02522_),
    .B1(_02524_),
    .B2(addr_i_3_),
    .Y(_02526_)
  );
  sg13g2_nor2_1 _12771_ (
    .A(_01612_),
    .B(_02526_),
    .Y(_02527_)
  );
  sg13g2_buf_1 _12772_ (
    .A(_09371_),
    .X(_02528_)
  );
  sg13g2_nand2_1 _12773_ (
    .A(_07933_),
    .B(_04937_),
    .Y(_02529_)
  );
  sg13g2_buf_1 _12774_ (
    .A(_01970_),
    .X(_02530_)
  );
  sg13g2_a21oi_1 _12775_ (
    .A1(_02528_),
    .A2(_02529_),
    .B1(_02530_),
    .Y(_02531_)
  );
  sg13g2_o21ai_1 _12776_ (
    .A1(_01582_),
    .A2(_02531_),
    .B1(addr_i_5_),
    .Y(_02532_)
  );
  sg13g2_nand2_1 _12777_ (
    .A(addr_i_5_),
    .B(_09393_),
    .Y(_02533_)
  );
  sg13g2_a21oi_1 _12778_ (
    .A1(_01240_),
    .A2(_02533_),
    .B1(_01660_),
    .Y(_02534_)
  );
  sg13g2_nand2_1 _12779_ (
    .A(addr_i_7_),
    .B(_00422_),
    .Y(_02535_)
  );
  sg13g2_a21oi_1 _12780_ (
    .A1(_02532_),
    .A2(_02534_),
    .B1(_02535_),
    .Y(_02537_)
  );
  sg13g2_a22oi_1 _12781_ (
    .A1(_02520_),
    .A2(_02527_),
    .B1(addr_i_12_),
    .B2(_02537_),
    .Y(_02538_)
  );
  sg13g2_nor2_1 _12782_ (
    .A(addr_i_9_),
    .B(_01760_),
    .Y(_02539_)
  );
  sg13g2_o21ai_1 _12783_ (
    .A1(_00158_),
    .A2(_09348_),
    .B1(_01528_),
    .Y(_02540_)
  );
  sg13g2_a21oi_1 _12784_ (
    .A1(_00339_),
    .A2(_02540_),
    .B1(_07149_),
    .Y(_02541_)
  );
  sg13g2_nor2_1 _12785_ (
    .A(_06840_),
    .B(_06485_),
    .Y(_02542_)
  );
  sg13g2_o21ai_1 _12786_ (
    .A1(_01112_),
    .A2(_02542_),
    .B1(_00485_),
    .Y(_02543_)
  );
  sg13g2_nand2_1 _12787_ (
    .A(_02048_),
    .B(_02543_),
    .Y(_02544_)
  );
  sg13g2_o21ai_1 _12788_ (
    .A1(_02541_),
    .A2(_02544_),
    .B1(_01119_),
    .Y(_02545_)
  );
  sg13g2_nand2_1 _12789_ (
    .A(_05281_),
    .B(_09050_),
    .Y(_02546_)
  );
  sg13g2_o21ai_1 _12790_ (
    .A1(_02076_),
    .A2(_07038_),
    .B1(_02546_),
    .Y(_02548_)
  );
  sg13g2_nand3_1 _12791_ (
    .A(addr_i_6_),
    .B(_03776_),
    .C(_01672_),
    .Y(_02549_)
  );
  sg13g2_a21oi_1 _12792_ (
    .A1(_01212_),
    .A2(_02549_),
    .B1(addr_i_3_),
    .Y(_02550_)
  );
  sg13g2_a22oi_1 _12793_ (
    .A1(addr_i_5_),
    .A2(_02548_),
    .B1(_02550_),
    .B2(_01194_),
    .Y(_02551_)
  );
  sg13g2_nand2_1 _12794_ (
    .A(addr_i_7_),
    .B(_01339_),
    .Y(_02552_)
  );
  sg13g2_nand3_1 _12795_ (
    .A(addr_i_3_),
    .B(_00199_),
    .C(_04804_),
    .Y(_02553_)
  );
  sg13g2_nand3_1 _12796_ (
    .A(addr_i_4_),
    .B(_00065_),
    .C(_03953_),
    .Y(_02554_)
  );
  sg13g2_a21oi_1 _12797_ (
    .A1(_02553_),
    .A2(_02554_),
    .B1(addr_i_6_),
    .Y(_02555_)
  );
  sg13g2_a22oi_1 _12798_ (
    .A1(_00192_),
    .A2(_02552_),
    .B1(_02555_),
    .B2(addr_i_8_),
    .Y(_02556_)
  );
  sg13g2_o21ai_1 _12799_ (
    .A1(addr_i_4_),
    .A2(_02551_),
    .B1(_02556_),
    .Y(_02557_)
  );
  sg13g2_a21oi_1 _12800_ (
    .A1(addr_i_2_),
    .A2(_02342_),
    .B1(_00559_),
    .Y(_02559_)
  );
  sg13g2_nand2_1 _12801_ (
    .A(addr_i_4_),
    .B(_00725_),
    .Y(_02560_)
  );
  sg13g2_nor2_1 _12802_ (
    .A(addr_i_3_),
    .B(_02268_),
    .Y(_02561_)
  );
  sg13g2_nand2_1 _12803_ (
    .A(_01310_),
    .B(_00353_),
    .Y(_02562_)
  );
  sg13g2_a21oi_1 _12804_ (
    .A1(_02560_),
    .A2(_02561_),
    .B1(_02562_),
    .Y(_02563_)
  );
  sg13g2_o21ai_1 _12805_ (
    .A1(_05877_),
    .A2(_02559_),
    .B1(_02563_),
    .Y(_02564_)
  );
  sg13g2_nand4_1 _12806_ (
    .A(addr_i_9_),
    .B(_02545_),
    .C(_02557_),
    .D(_02564_),
    .Y(_02565_)
  );
  sg13g2_nand2b_1 _12807_ (
    .A_N(_02539_),
    .B(_02565_),
    .Y(_02566_)
  );
  sg13g2_nand2_1 _12808_ (
    .A(_01527_),
    .B(_09415_),
    .Y(_02567_)
  );
  sg13g2_a22oi_1 _12809_ (
    .A1(addr_i_4_),
    .A2(_02567_),
    .B1(_00426_),
    .B2(_01380_),
    .Y(_02568_)
  );
  sg13g2_a21oi_1 _12810_ (
    .A1(_01815_),
    .A2(_02187_),
    .B1(_00726_),
    .Y(_02570_)
  );
  sg13g2_a22oi_1 _12811_ (
    .A1(addr_i_6_),
    .A2(_02560_),
    .B1(_02570_),
    .B2(_03227_),
    .Y(_02571_)
  );
  sg13g2_o21ai_1 _12812_ (
    .A1(addr_i_3_),
    .A2(_02568_),
    .B1(_02571_),
    .Y(_02572_)
  );
  sg13g2_nand2_1 _12813_ (
    .A(addr_i_3_),
    .B(_05025_),
    .Y(_02573_)
  );
  sg13g2_o21ai_1 _12814_ (
    .A1(_00454_),
    .A2(_04119_),
    .B1(_00648_),
    .Y(_02574_)
  );
  sg13g2_a21o_1 _12815_ (
    .A1(_02573_),
    .A2(_02574_),
    .B1(addr_i_6_),
    .X(_02575_)
  );
  sg13g2_a21oi_1 _12816_ (
    .A1(_00298_),
    .A2(_01232_),
    .B1(addr_i_8_),
    .Y(_02576_)
  );
  sg13g2_buf_1 _12817_ (
    .A(_00679_),
    .X(_02577_)
  );
  sg13g2_buf_1 _12818_ (
    .A(_00543_),
    .X(_02578_)
  );
  sg13g2_nand4_1 _12819_ (
    .A(_00505_),
    .B(_02577_),
    .C(_00080_),
    .D(_02578_),
    .Y(_02579_)
  );
  sg13g2_o21ai_1 _12820_ (
    .A1(_00132_),
    .A2(_01246_),
    .B1(addr_i_5_),
    .Y(_02581_)
  );
  sg13g2_nand4_1 _12821_ (
    .A(_02575_),
    .B(_02576_),
    .C(_02579_),
    .D(_02581_),
    .Y(_02582_)
  );
  sg13g2_nand2_1 _12822_ (
    .A(addr_i_5_),
    .B(_03743_),
    .Y(_02583_)
  );
  sg13g2_nor2_1 _12823_ (
    .A(_02191_),
    .B(_02583_),
    .Y(_02584_)
  );
  sg13g2_o21ai_1 _12824_ (
    .A1(_04550_),
    .A2(_03490_),
    .B1(_04075_),
    .Y(_02585_)
  );
  sg13g2_nor2_1 _12825_ (
    .A(_08343_),
    .B(_00578_),
    .Y(_02586_)
  );
  sg13g2_a21oi_1 _12826_ (
    .A1(addr_i_4_),
    .A2(_02585_),
    .B1(_02586_),
    .Y(_02587_)
  );
  sg13g2_nor2_1 _12827_ (
    .A(addr_i_3_),
    .B(_02587_),
    .Y(_02588_)
  );
  sg13g2_o21ai_1 _12828_ (
    .A1(_02584_),
    .A2(_02588_),
    .B1(_01118_),
    .Y(_02589_)
  );
  sg13g2_nand3_1 _12829_ (
    .A(_02572_),
    .B(_02582_),
    .C(_02589_),
    .Y(_02590_)
  );
  sg13g2_nor2_1 _12830_ (
    .A(addr_i_6_),
    .B(_01228_),
    .Y(_02592_)
  );
  sg13g2_a21o_1 _12831_ (
    .A1(addr_i_3_),
    .A2(_02592_),
    .B1(_02215_),
    .X(_02593_)
  );
  sg13g2_a21oi_1 _12832_ (
    .A1(_06884_),
    .A2(_02369_),
    .B1(_09506_),
    .Y(_02594_)
  );
  sg13g2_o21ai_1 _12833_ (
    .A1(addr_i_2_),
    .A2(_01585_),
    .B1(_01653_),
    .Y(_02595_)
  );
  sg13g2_o21ai_1 _12834_ (
    .A1(addr_i_2_),
    .A2(_02594_),
    .B1(_02595_),
    .Y(_02596_)
  );
  sg13g2_o21ai_1 _12835_ (
    .A1(_08188_),
    .A2(_01015_),
    .B1(_00607_),
    .Y(_02597_)
  );
  sg13g2_buf_1 _12836_ (
    .A(_00742_),
    .X(_02598_)
  );
  sg13g2_o21ai_1 _12837_ (
    .A1(_02598_),
    .A2(_06574_),
    .B1(addr_i_7_),
    .Y(_02599_)
  );
  sg13g2_a21oi_1 _12838_ (
    .A1(_02597_),
    .A2(_02599_),
    .B1(addr_i_4_),
    .Y(_02600_)
  );
  sg13g2_a221oi_1 _12839_ (
    .A1(addr_i_2_),
    .A2(_02593_),
    .B1(_02596_),
    .B2(addr_i_4_),
    .C1(_02600_),
    .Y(_02601_)
  );
  sg13g2_o21ai_1 _12840_ (
    .A1(_00703_),
    .A2(_00051_),
    .B1(_02601_),
    .Y(_02603_)
  );
  sg13g2_buf_1 _12841_ (
    .A(_02952_),
    .X(_02604_)
  );
  sg13g2_a22oi_1 _12842_ (
    .A1(_07149_),
    .A2(_00409_),
    .B1(_00214_),
    .B2(_00230_),
    .Y(_02605_)
  );
  sg13g2_nand2_1 _12843_ (
    .A(_02165_),
    .B(_02605_),
    .Y(_02606_)
  );
  sg13g2_nor2_1 _12844_ (
    .A(addr_i_7_),
    .B(_00213_),
    .Y(_02607_)
  );
  sg13g2_nand3_1 _12845_ (
    .A(_01616_),
    .B(_01464_),
    .C(_02607_),
    .Y(_02608_)
  );
  sg13g2_a21oi_1 _12846_ (
    .A1(addr_i_3_),
    .A2(_00477_),
    .B1(_00322_),
    .Y(_02609_)
  );
  sg13g2_a21oi_1 _12847_ (
    .A1(_06806_),
    .A2(_00712_),
    .B1(_02171_),
    .Y(_02610_)
  );
  sg13g2_o21ai_1 _12848_ (
    .A1(_02277_),
    .A2(_02609_),
    .B1(_02610_),
    .Y(_02611_)
  );
  sg13g2_nand3_1 _12849_ (
    .A(addr_i_5_),
    .B(_01518_),
    .C(_02611_),
    .Y(_02612_)
  );
  sg13g2_nand4_1 _12850_ (
    .A(addr_i_12_),
    .B(_02606_),
    .C(_02608_),
    .D(_02612_),
    .Y(_02614_)
  );
  sg13g2_a221oi_1 _12851_ (
    .A1(addr_i_9_),
    .A2(_02590_),
    .B1(_02603_),
    .B2(_02604_),
    .C1(_02614_),
    .Y(_02615_)
  );
  sg13g2_a22oi_1 _12852_ (
    .A1(_02538_),
    .A2(_02566_),
    .B1(_02615_),
    .B2(addr_i_10_),
    .Y(_02616_)
  );
  sg13g2_a22oi_1 _12853_ (
    .A1(addr_i_10_),
    .A2(_02512_),
    .B1(_02616_),
    .B2(addr_i_11_),
    .Y(_02617_)
  );
  sg13g2_a21oi_1 _12854_ (
    .A1(_02365_),
    .A2(_02402_),
    .B1(_02617_),
    .Y(data_o_15_)
  );
  sg13g2_nand2_1 _12855_ (
    .A(_06972_),
    .B(_01004_),
    .Y(_02618_)
  );
  sg13g2_a21oi_1 _12856_ (
    .A1(addr_i_6_),
    .A2(_04494_),
    .B1(addr_i_2_),
    .Y(_02619_)
  );
  sg13g2_a21oi_1 _12857_ (
    .A1(_00316_),
    .A2(_05457_),
    .B1(_08696_),
    .Y(_02620_)
  );
  sg13g2_a22oi_1 _12858_ (
    .A1(addr_i_4_),
    .A2(_02618_),
    .B1(_02619_),
    .B2(_02620_),
    .Y(_02621_)
  );
  sg13g2_nor2_1 _12859_ (
    .A(_02371_),
    .B(_02733_),
    .Y(_02622_)
  );
  sg13g2_o21ai_1 _12860_ (
    .A1(_00072_),
    .A2(_02622_),
    .B1(addr_i_6_),
    .Y(_02624_)
  );
  sg13g2_o21ai_1 _12861_ (
    .A1(_05867_),
    .A2(_02621_),
    .B1(_02624_),
    .Y(_02625_)
  );
  sg13g2_nor2_1 _12862_ (
    .A(_07491_),
    .B(_02108_),
    .Y(_02626_)
  );
  sg13g2_nor2_1 _12863_ (
    .A(_00165_),
    .B(_02626_),
    .Y(_02627_)
  );
  sg13g2_o21ai_1 _12864_ (
    .A1(addr_i_3_),
    .A2(_02627_),
    .B1(_00056_),
    .Y(_02628_)
  );
  sg13g2_nand3_1 _12865_ (
    .A(addr_i_4_),
    .B(_00994_),
    .C(_01230_),
    .Y(_02629_)
  );
  sg13g2_o21ai_1 _12866_ (
    .A1(addr_i_4_),
    .A2(_02628_),
    .B1(_02629_),
    .Y(_02630_)
  );
  sg13g2_nand2b_1 _12867_ (
    .A_N(_02625_),
    .B(_02630_),
    .Y(_02631_)
  );
  sg13g2_nor2_1 _12868_ (
    .A(_00044_),
    .B(_02558_),
    .Y(_02632_)
  );
  sg13g2_nor2_1 _12869_ (
    .A(_05070_),
    .B(_08531_),
    .Y(_02633_)
  );
  sg13g2_o21ai_1 _12870_ (
    .A1(_02632_),
    .A2(_02633_),
    .B1(addr_i_3_),
    .Y(_02635_)
  );
  sg13g2_o21ai_1 _12871_ (
    .A1(_08266_),
    .A2(_09504_),
    .B1(_02635_),
    .Y(_02636_)
  );
  sg13g2_o21ai_1 _12872_ (
    .A1(_00380_),
    .A2(_00025_),
    .B1(_04384_),
    .Y(_02637_)
  );
  sg13g2_nor2_1 _12873_ (
    .A(_00199_),
    .B(_00099_),
    .Y(_02638_)
  );
  sg13g2_nor3_1 _12874_ (
    .A(addr_i_4_),
    .B(addr_i_7_),
    .C(addr_i_6_),
    .Y(_02639_)
  );
  sg13g2_a221oi_1 _12875_ (
    .A1(addr_i_3_),
    .A2(_02637_),
    .B1(_02638_),
    .B2(_00616_),
    .C1(_02639_),
    .Y(_02640_)
  );
  sg13g2_nor2_1 _12876_ (
    .A(_05700_),
    .B(_07160_),
    .Y(_02641_)
  );
  sg13g2_o21ai_1 _12877_ (
    .A1(_00010_),
    .A2(_02641_),
    .B1(_00268_),
    .Y(_02642_)
  );
  sg13g2_o21ai_1 _12878_ (
    .A1(addr_i_2_),
    .A2(_02640_),
    .B1(_02642_),
    .Y(_02643_)
  );
  sg13g2_a22oi_1 _12879_ (
    .A1(addr_i_2_),
    .A2(_02636_),
    .B1(_02643_),
    .B2(addr_i_8_),
    .Y(_02644_)
  );
  sg13g2_a21o_1 _12880_ (
    .A1(addr_i_8_),
    .A2(_02631_),
    .B1(_02644_),
    .X(_02646_)
  );
  sg13g2_o21ai_1 _12881_ (
    .A1(addr_i_2_),
    .A2(_09050_),
    .B1(addr_i_5_),
    .Y(_02647_)
  );
  sg13g2_a21oi_1 _12882_ (
    .A1(_01077_),
    .A2(_02647_),
    .B1(addr_i_3_),
    .Y(_02648_)
  );
  sg13g2_a21oi_1 _12883_ (
    .A1(_07779_),
    .A2(_02218_),
    .B1(addr_i_2_),
    .Y(_02649_)
  );
  sg13g2_a21oi_1 _12884_ (
    .A1(_00050_),
    .A2(_01441_),
    .B1(_00046_),
    .Y(_02650_)
  );
  sg13g2_nor4_1 _12885_ (
    .A(_09498_),
    .B(_02648_),
    .C(_02649_),
    .D(_02650_),
    .Y(_02651_)
  );
  sg13g2_nor3_1 _12886_ (
    .A(addr_i_3_),
    .B(addr_i_7_),
    .C(addr_i_6_),
    .Y(_02652_)
  );
  sg13g2_nor3_1 _12887_ (
    .A(_00535_),
    .B(_06729_),
    .C(_07105_),
    .Y(_02653_)
  );
  sg13g2_o21ai_1 _12888_ (
    .A1(_02652_),
    .A2(_02653_),
    .B1(addr_i_5_),
    .Y(_02654_)
  );
  sg13g2_o21ai_1 _12889_ (
    .A1(_01194_),
    .A2(_01711_),
    .B1(addr_i_6_),
    .Y(_02655_)
  );
  sg13g2_a21oi_1 _12890_ (
    .A1(_02654_),
    .A2(_02655_),
    .B1(addr_i_4_),
    .Y(_02657_)
  );
  sg13g2_a21o_1 _12891_ (
    .A1(addr_i_4_),
    .A2(_02651_),
    .B1(_02657_),
    .X(_02658_)
  );
  sg13g2_nand2_1 _12892_ (
    .A(_00899_),
    .B(_01499_),
    .Y(_02659_)
  );
  sg13g2_nand2_1 _12893_ (
    .A(_06695_),
    .B(_00131_),
    .Y(_02660_)
  );
  sg13g2_nand2_1 _12894_ (
    .A(_05524_),
    .B(_09485_),
    .Y(_02661_)
  );
  sg13g2_o21ai_1 _12895_ (
    .A1(_01086_),
    .A2(_00132_),
    .B1(addr_i_5_),
    .Y(_02662_)
  );
  sg13g2_a21oi_1 _12896_ (
    .A1(_02661_),
    .A2(_02662_),
    .B1(_01935_),
    .Y(_02663_)
  );
  sg13g2_a22oi_1 _12897_ (
    .A1(addr_i_2_),
    .A2(_02659_),
    .B1(_02660_),
    .B2(_02663_),
    .Y(_02664_)
  );
  sg13g2_o21ai_1 _12898_ (
    .A1(_00492_),
    .A2(_07558_),
    .B1(_00249_),
    .Y(_02665_)
  );
  sg13g2_nand2_1 _12899_ (
    .A(addr_i_7_),
    .B(_02472_),
    .Y(_02666_)
  );
  sg13g2_a21oi_1 _12900_ (
    .A1(_01386_),
    .A2(_02666_),
    .B1(addr_i_3_),
    .Y(_02668_)
  );
  sg13g2_o21ai_1 _12901_ (
    .A1(_02665_),
    .A2(_02668_),
    .B1(_01324_),
    .Y(_02669_)
  );
  sg13g2_a221oi_1 _12902_ (
    .A1(addr_i_8_),
    .A2(_02658_),
    .B1(_02664_),
    .B2(_02669_),
    .C1(addr_i_9_),
    .Y(_02670_)
  );
  sg13g2_a21o_1 _12903_ (
    .A1(addr_i_9_),
    .A2(_02646_),
    .B1(_02670_),
    .X(_02671_)
  );
  sg13g2_nand2_1 _12904_ (
    .A(addr_i_5_),
    .B(_00447_),
    .Y(_02672_)
  );
  sg13g2_nor2_1 _12905_ (
    .A(addr_i_3_),
    .B(_02672_),
    .Y(_02673_)
  );
  sg13g2_a22oi_1 _12906_ (
    .A1(addr_i_3_),
    .A2(_01164_),
    .B1(_02673_),
    .B2(_01837_),
    .Y(_02674_)
  );
  sg13g2_nand2_1 _12907_ (
    .A(_04461_),
    .B(_00687_),
    .Y(_02675_)
  );
  sg13g2_a21oi_1 _12908_ (
    .A1(_00401_),
    .A2(_02675_),
    .B1(_01082_),
    .Y(_02676_)
  );
  sg13g2_o21ai_1 _12909_ (
    .A1(_01630_),
    .A2(_02674_),
    .B1(_02676_),
    .Y(_02677_)
  );
  sg13g2_a21oi_1 _12910_ (
    .A1(_02755_),
    .A2(_01355_),
    .B1(_01041_),
    .Y(_02679_)
  );
  sg13g2_nand3_1 _12911_ (
    .A(_00314_),
    .B(_02498_),
    .C(_02679_),
    .Y(_02680_)
  );
  sg13g2_nand3_1 _12912_ (
    .A(_02501_),
    .B(_01453_),
    .C(_00852_),
    .Y(_02681_)
  );
  sg13g2_nand3_1 _12913_ (
    .A(addr_i_9_),
    .B(_02680_),
    .C(_02681_),
    .Y(_02682_)
  );
  sg13g2_nand2_1 _12914_ (
    .A(addr_i_4_),
    .B(_04937_),
    .Y(_02683_)
  );
  sg13g2_nand2_1 _12915_ (
    .A(_00371_),
    .B(_02683_),
    .Y(_02684_)
  );
  sg13g2_nor2_1 _12916_ (
    .A(addr_i_2_),
    .B(_00008_),
    .Y(_02685_)
  );
  sg13g2_nand2_1 _12917_ (
    .A(_01169_),
    .B(_02685_),
    .Y(_02686_)
  );
  sg13g2_a21oi_1 _12918_ (
    .A1(_00339_),
    .A2(_02686_),
    .B1(addr_i_6_),
    .Y(_02687_)
  );
  sg13g2_a22oi_1 _12919_ (
    .A1(addr_i_3_),
    .A2(_02684_),
    .B1(_02687_),
    .B2(_03062_),
    .Y(_02688_)
  );
  sg13g2_nand3_1 _12920_ (
    .A(addr_i_3_),
    .B(addr_i_4_),
    .C(_08774_),
    .Y(_02690_)
  );
  sg13g2_o21ai_1 _12921_ (
    .A1(addr_i_4_),
    .A2(_01555_),
    .B1(_02690_),
    .Y(_02691_)
  );
  sg13g2_a22oi_1 _12922_ (
    .A1(_01324_),
    .A2(_02691_),
    .B1(_00885_),
    .B2(_01391_),
    .Y(_02692_)
  );
  sg13g2_nor3_1 _12923_ (
    .A(_02682_),
    .B(_02688_),
    .C(_02692_),
    .Y(_02693_)
  );
  sg13g2_buf_1 _12924_ (
    .A(_01175_),
    .X(_02694_)
  );
  sg13g2_nand2_1 _12925_ (
    .A(_02152_),
    .B(_03194_),
    .Y(_02695_)
  );
  sg13g2_o21ai_1 _12926_ (
    .A1(_08896_),
    .A2(_03172_),
    .B1(_08044_),
    .Y(_02696_)
  );
  sg13g2_nand3_1 _12927_ (
    .A(_02694_),
    .B(_02695_),
    .C(_02696_),
    .Y(_02697_)
  );
  sg13g2_nor2_1 _12928_ (
    .A(_06884_),
    .B(_00543_),
    .Y(_02698_)
  );
  sg13g2_a22oi_1 _12929_ (
    .A1(addr_i_3_),
    .A2(_02697_),
    .B1(_02698_),
    .B2(_01391_),
    .Y(_02699_)
  );
  sg13g2_o21ai_1 _12930_ (
    .A1(_01024_),
    .A2(_02203_),
    .B1(addr_i_3_),
    .Y(_02701_)
  );
  sg13g2_o21ai_1 _12931_ (
    .A1(addr_i_4_),
    .A2(_00223_),
    .B1(_00022_),
    .Y(_02702_)
  );
  sg13g2_nand3_1 _12932_ (
    .A(_01425_),
    .B(_02701_),
    .C(_02702_),
    .Y(_02703_)
  );
  sg13g2_o21ai_1 _12933_ (
    .A1(_03238_),
    .A2(_02703_),
    .B1(_00396_),
    .Y(_02704_)
  );
  sg13g2_a22oi_1 _12934_ (
    .A1(addr_i_2_),
    .A2(_08553_),
    .B1(_06010_),
    .B2(addr_i_3_),
    .Y(_02705_)
  );
  sg13g2_a22oi_1 _12935_ (
    .A1(addr_i_4_),
    .A2(_00993_),
    .B1(_01049_),
    .B2(_01935_),
    .Y(_02706_)
  );
  sg13g2_o21ai_1 _12936_ (
    .A1(_02705_),
    .A2(_02706_),
    .B1(_00610_),
    .Y(_02707_)
  );
  sg13g2_nand2_1 _12937_ (
    .A(addr_i_3_),
    .B(_00303_),
    .Y(_02708_)
  );
  sg13g2_o21ai_1 _12938_ (
    .A1(addr_i_4_),
    .A2(_02514_),
    .B1(_01277_),
    .Y(_02709_)
  );
  sg13g2_nand4_1 _12939_ (
    .A(_09105_),
    .B(_02708_),
    .C(_01182_),
    .D(_02709_),
    .Y(_02710_)
  );
  sg13g2_o21ai_1 _12940_ (
    .A1(_02261_),
    .A2(_02710_),
    .B1(_00440_),
    .Y(_02712_)
  );
  sg13g2_nand2_1 _12941_ (
    .A(_02707_),
    .B(_02712_),
    .Y(_02713_)
  );
  sg13g2_nor3_1 _12942_ (
    .A(_02699_),
    .B(_02704_),
    .C(_02713_),
    .Y(_02714_)
  );
  sg13g2_a22oi_1 _12943_ (
    .A1(_02677_),
    .A2(_02693_),
    .B1(_02714_),
    .B2(addr_i_10_),
    .Y(_02715_)
  );
  sg13g2_a22oi_1 _12944_ (
    .A1(addr_i_10_),
    .A2(_02671_),
    .B1(_02715_),
    .B2(addr_i_11_),
    .Y(_02716_)
  );
  sg13g2_nor3_1 _12945_ (
    .A(_00243_),
    .B(addr_i_5_),
    .C(_01861_),
    .Y(_02717_)
  );
  sg13g2_inv_1 _12946_ (
    .A(_01374_),
    .Y(_02718_)
  );
  sg13g2_nand2_1 _12947_ (
    .A(_00228_),
    .B(_02930_),
    .Y(_02719_)
  );
  sg13g2_nand3_1 _12948_ (
    .A(addr_i_2_),
    .B(_00147_),
    .C(_03325_),
    .Y(_02720_)
  );
  sg13g2_a21oi_1 _12949_ (
    .A1(_00185_),
    .A2(_02720_),
    .B1(_00485_),
    .Y(_02721_)
  );
  sg13g2_a22oi_1 _12950_ (
    .A1(_07149_),
    .A2(_02719_),
    .B1(_02721_),
    .B2(_07425_),
    .Y(_02723_)
  );
  sg13g2_nor2_1 _12951_ (
    .A(_00290_),
    .B(_02723_),
    .Y(_02724_)
  );
  sg13g2_nand2_1 _12952_ (
    .A(_00956_),
    .B(_03545_),
    .Y(_02725_)
  );
  sg13g2_nand2_1 _12953_ (
    .A(_00353_),
    .B(_02725_),
    .Y(_02726_)
  );
  sg13g2_o21ai_1 _12954_ (
    .A1(_00491_),
    .A2(_05125_),
    .B1(addr_i_4_),
    .Y(_02727_)
  );
  sg13g2_a22oi_1 _12955_ (
    .A1(addr_i_10_),
    .A2(_06375_),
    .B1(_00791_),
    .B2(_02268_),
    .Y(_02728_)
  );
  sg13g2_nand2_1 _12956_ (
    .A(_02727_),
    .B(_02728_),
    .Y(_02729_)
  );
  sg13g2_a21oi_1 _12957_ (
    .A1(addr_i_3_),
    .A2(_02726_),
    .B1(_02729_),
    .Y(_02730_)
  );
  sg13g2_a21oi_1 _12958_ (
    .A1(_06132_),
    .A2(_00785_),
    .B1(_00700_),
    .Y(_02731_)
  );
  sg13g2_buf_1 _12959_ (
    .A(_06884_),
    .X(_02732_)
  );
  sg13g2_nor2_1 _12960_ (
    .A(_00467_),
    .B(_02732_),
    .Y(_02734_)
  );
  sg13g2_nor2_1 _12961_ (
    .A(_02731_),
    .B(_02734_),
    .Y(_02735_)
  );
  sg13g2_nor2_1 _12962_ (
    .A(_01034_),
    .B(_02735_),
    .Y(_02736_)
  );
  sg13g2_nor4_1 _12963_ (
    .A(_02718_),
    .B(_02724_),
    .C(_02730_),
    .D(_02736_),
    .Y(_02737_)
  );
  sg13g2_nand2_1 _12964_ (
    .A(_00840_),
    .B(_09061_),
    .Y(_02738_)
  );
  sg13g2_o21ai_1 _12965_ (
    .A1(_01355_),
    .A2(_02738_),
    .B1(addr_i_10_),
    .Y(_02739_)
  );
  sg13g2_o21ai_1 _12966_ (
    .A1(_02717_),
    .A2(_02737_),
    .B1(_02739_),
    .Y(_02740_)
  );
  sg13g2_a21o_1 _12967_ (
    .A1(addr_i_11_),
    .A2(_02740_),
    .B1(_00812_),
    .X(_02741_)
  );
  sg13g2_buf_1 _12968_ (
    .A(_01954_),
    .X(_02742_)
  );
  sg13g2_o21ai_1 _12969_ (
    .A1(_01500_),
    .A2(_01754_),
    .B1(_02742_),
    .Y(_02743_)
  );
  sg13g2_nand2_1 _12970_ (
    .A(_00440_),
    .B(_02743_),
    .Y(_02745_)
  );
  sg13g2_nand2_1 _12971_ (
    .A(addr_i_4_),
    .B(_00711_),
    .Y(_02746_)
  );
  sg13g2_a21oi_1 _12972_ (
    .A1(_02467_),
    .A2(_02746_),
    .B1(addr_i_5_),
    .Y(_02747_)
  );
  sg13g2_o21ai_1 _12973_ (
    .A1(_02441_),
    .A2(_00177_),
    .B1(addr_i_3_),
    .Y(_02748_)
  );
  sg13g2_o21ai_1 _12974_ (
    .A1(addr_i_2_),
    .A2(_01019_),
    .B1(_07547_),
    .Y(_02749_)
  );
  sg13g2_nor2_1 _12975_ (
    .A(addr_i_6_),
    .B(_00252_),
    .Y(_02750_)
  );
  sg13g2_o21ai_1 _12976_ (
    .A1(addr_i_3_),
    .A2(_02750_),
    .B1(_00695_),
    .Y(_02751_)
  );
  sg13g2_nand2_1 _12977_ (
    .A(_00497_),
    .B(_02751_),
    .Y(_02752_)
  );
  sg13g2_nand4_1 _12978_ (
    .A(_00610_),
    .B(_02748_),
    .C(_02749_),
    .D(_02752_),
    .Y(_02753_)
  );
  sg13g2_o21ai_1 _12979_ (
    .A1(_02745_),
    .A2(_02747_),
    .B1(_02753_),
    .Y(_02754_)
  );
  sg13g2_a21oi_1 _12980_ (
    .A1(_02136_),
    .A2(_07094_),
    .B1(addr_i_5_),
    .Y(_02756_)
  );
  sg13g2_o21ai_1 _12981_ (
    .A1(_03150_),
    .A2(_02756_),
    .B1(addr_i_2_),
    .Y(_02757_)
  );
  sg13g2_nand2_1 _12982_ (
    .A(_01410_),
    .B(_02757_),
    .Y(_02758_)
  );
  sg13g2_buf_1 _12983_ (
    .A(_00006_),
    .X(_02759_)
  );
  sg13g2_a22oi_1 _12984_ (
    .A1(_00015_),
    .A2(_02759_),
    .B1(_01542_),
    .B2(_01520_),
    .Y(_02760_)
  );
  sg13g2_nand2_1 _12985_ (
    .A(_02053_),
    .B(_06077_),
    .Y(_02761_)
  );
  sg13g2_a21oi_1 _12986_ (
    .A1(addr_i_2_),
    .A2(_02761_),
    .B1(addr_i_4_),
    .Y(_02762_)
  );
  sg13g2_nor3_1 _12987_ (
    .A(addr_i_3_),
    .B(_02760_),
    .C(_02762_),
    .Y(_02763_)
  );
  sg13g2_o21ai_1 _12988_ (
    .A1(_00930_),
    .A2(_08553_),
    .B1(addr_i_8_),
    .Y(_02764_)
  );
  sg13g2_a22oi_1 _12989_ (
    .A1(addr_i_3_),
    .A2(_02758_),
    .B1(_02763_),
    .B2(_02764_),
    .Y(_02765_)
  );
  sg13g2_o21ai_1 _12990_ (
    .A1(_02754_),
    .A2(_02765_),
    .B1(_05214_),
    .Y(_02767_)
  );
  sg13g2_o21ai_1 _12991_ (
    .A1(_00515_),
    .A2(_01787_),
    .B1(addr_i_2_),
    .Y(_02768_)
  );
  sg13g2_a22oi_1 _12992_ (
    .A1(addr_i_4_),
    .A2(_00328_),
    .B1(_02203_),
    .B2(_07425_),
    .Y(_02769_)
  );
  sg13g2_nand2b_1 _12993_ (
    .A_N(_02769_),
    .B(addr_i_3_),
    .Y(_02770_)
  );
  sg13g2_nand4_1 _12994_ (
    .A(_00708_),
    .B(_00907_),
    .C(_02768_),
    .D(_02770_),
    .Y(_02771_)
  );
  sg13g2_buf_1 _12995_ (
    .A(_08288_),
    .X(_02772_)
  );
  sg13g2_o21ai_1 _12996_ (
    .A1(_02772_),
    .A2(_00885_),
    .B1(addr_i_4_),
    .Y(_02773_)
  );
  sg13g2_nor2_1 _12997_ (
    .A(addr_i_4_),
    .B(_00591_),
    .Y(_02774_)
  );
  sg13g2_a21oi_1 _12998_ (
    .A1(addr_i_3_),
    .A2(_02774_),
    .B1(_00588_),
    .Y(_02775_)
  );
  sg13g2_o21ai_1 _12999_ (
    .A1(_02261_),
    .A2(_01986_),
    .B1(_04052_),
    .Y(_02776_)
  );
  sg13g2_nand3_1 _13000_ (
    .A(_02773_),
    .B(_02775_),
    .C(_02776_),
    .Y(_02778_)
  );
  sg13g2_a22oi_1 _13001_ (
    .A1(addr_i_4_),
    .A2(_02382_),
    .B1(_01560_),
    .B2(_01282_),
    .Y(_02779_)
  );
  sg13g2_nand2b_1 _13002_ (
    .A_N(addr_i_8_),
    .B(addr_i_6_),
    .Y(_02780_)
  );
  sg13g2_buf_1 _13003_ (
    .A(_02780_),
    .X(_02781_)
  );
  sg13g2_nor3_1 _13004_ (
    .A(_05833_),
    .B(_02781_),
    .C(_02622_),
    .Y(_02782_)
  );
  sg13g2_o21ai_1 _13005_ (
    .A1(addr_i_3_),
    .A2(_02779_),
    .B1(_02782_),
    .Y(_02783_)
  );
  sg13g2_o21ai_1 _13006_ (
    .A1(_07879_),
    .A2(_06010_),
    .B1(addr_i_3_),
    .Y(_02784_)
  );
  sg13g2_nand2_1 _13007_ (
    .A(_06851_),
    .B(_00571_),
    .Y(_02785_)
  );
  sg13g2_a21oi_1 _13008_ (
    .A1(_00200_),
    .A2(_02785_),
    .B1(_01015_),
    .Y(_02786_)
  );
  sg13g2_nand2_1 _13009_ (
    .A(_02784_),
    .B(_02786_),
    .Y(_02787_)
  );
  sg13g2_a22oi_1 _13010_ (
    .A1(_06873_),
    .A2(_02490_),
    .B1(_05568_),
    .B2(_04672_),
    .Y(_02789_)
  );
  sg13g2_a22oi_1 _13011_ (
    .A1(_01633_),
    .A2(_02787_),
    .B1(_02789_),
    .B2(addr_i_9_),
    .Y(_02790_)
  );
  sg13g2_nand4_1 _13012_ (
    .A(_02771_),
    .B(_02778_),
    .C(_02783_),
    .D(_02790_),
    .Y(_02791_)
  );
  sg13g2_nor2_1 _13013_ (
    .A(addr_i_3_),
    .B(_08863_),
    .Y(_02792_)
  );
  sg13g2_o21ai_1 _13014_ (
    .A1(_01787_),
    .A2(_02792_),
    .B1(addr_i_2_),
    .Y(_02793_)
  );
  sg13g2_nor2_1 _13015_ (
    .A(_02471_),
    .B(_06032_),
    .Y(_02794_)
  );
  sg13g2_a22oi_1 _13016_ (
    .A1(_00727_),
    .A2(_02369_),
    .B1(_02794_),
    .B2(addr_i_6_),
    .Y(_02795_)
  );
  sg13g2_buf_1 _13017_ (
    .A(_04041_),
    .X(_02796_)
  );
  sg13g2_a21oi_1 _13018_ (
    .A1(_00186_),
    .A2(_00926_),
    .B1(addr_i_3_),
    .Y(_02797_)
  );
  sg13g2_nor3_1 _13019_ (
    .A(_02796_),
    .B(_01977_),
    .C(_02797_),
    .Y(_02798_)
  );
  sg13g2_a21oi_1 _13020_ (
    .A1(_02793_),
    .A2(_02795_),
    .B1(_02798_),
    .Y(_02800_)
  );
  sg13g2_nor2_1 _13021_ (
    .A(_04318_),
    .B(_02733_),
    .Y(_02801_)
  );
  sg13g2_nor2_1 _13022_ (
    .A(_08045_),
    .B(_02801_),
    .Y(_02802_)
  );
  sg13g2_buf_1 _13023_ (
    .A(_04373_),
    .X(_02803_)
  );
  sg13g2_nand2_1 _13024_ (
    .A(_00001_),
    .B(_08852_),
    .Y(_02804_)
  );
  sg13g2_nand3_1 _13025_ (
    .A(_00211_),
    .B(_01555_),
    .C(_02804_),
    .Y(_02805_)
  );
  sg13g2_nand2_1 _13026_ (
    .A(addr_i_8_),
    .B(_00358_),
    .Y(_02806_)
  );
  sg13g2_nand2_1 _13027_ (
    .A(_03380_),
    .B(_02141_),
    .Y(_02807_)
  );
  sg13g2_nor2_1 _13028_ (
    .A(_02053_),
    .B(_09493_),
    .Y(_02808_)
  );
  sg13g2_a221oi_1 _13029_ (
    .A1(_00731_),
    .A2(_01585_),
    .B1(_00010_),
    .B2(_02807_),
    .C1(_02808_),
    .Y(_02809_)
  );
  sg13g2_a22oi_1 _13030_ (
    .A1(_02803_),
    .A2(_02805_),
    .B1(_02806_),
    .B2(_02809_),
    .Y(_02811_)
  );
  sg13g2_a22oi_1 _13031_ (
    .A1(_02028_),
    .A2(_02802_),
    .B1(_02811_),
    .B2(_04705_),
    .Y(_02812_)
  );
  sg13g2_o21ai_1 _13032_ (
    .A1(addr_i_8_),
    .A2(_02800_),
    .B1(_02812_),
    .Y(_02813_)
  );
  sg13g2_nand3_1 _13033_ (
    .A(_00511_),
    .B(_02791_),
    .C(_02813_),
    .Y(_02814_)
  );
  sg13g2_buf_1 _13034_ (
    .A(_01757_),
    .X(_02815_)
  );
  sg13g2_a21oi_1 _13035_ (
    .A1(_02577_),
    .A2(_02815_),
    .B1(_00726_),
    .Y(_02816_)
  );
  sg13g2_o21ai_1 _13036_ (
    .A1(_00474_),
    .A2(_02816_),
    .B1(addr_i_4_),
    .Y(_02817_)
  );
  sg13g2_nand3_1 _13037_ (
    .A(_02803_),
    .B(_00351_),
    .C(_00140_),
    .Y(_02818_)
  );
  sg13g2_a21oi_1 _13038_ (
    .A1(_02817_),
    .A2(_02818_),
    .B1(addr_i_2_),
    .Y(_02819_)
  );
  sg13g2_nand2_1 _13039_ (
    .A(addr_i_5_),
    .B(_01309_),
    .Y(_02820_)
  );
  sg13g2_nand2_1 _13040_ (
    .A(_04362_),
    .B(_00154_),
    .Y(_02822_)
  );
  sg13g2_o21ai_1 _13041_ (
    .A1(_00183_),
    .A2(_01888_),
    .B1(_02514_),
    .Y(_02823_)
  );
  sg13g2_nand2_1 _13042_ (
    .A(_02822_),
    .B(_02823_),
    .Y(_02824_)
  );
  sg13g2_o21ai_1 _13043_ (
    .A1(addr_i_5_),
    .A2(_00183_),
    .B1(addr_i_2_),
    .Y(_02825_)
  );
  sg13g2_a21oi_1 _13044_ (
    .A1(_02577_),
    .A2(_02825_),
    .B1(addr_i_3_),
    .Y(_02826_)
  );
  sg13g2_o21ai_1 _13045_ (
    .A1(_02824_),
    .A2(_02826_),
    .B1(_00388_),
    .Y(_02827_)
  );
  sg13g2_o21ai_1 _13046_ (
    .A1(_00103_),
    .A2(_02820_),
    .B1(_02827_),
    .Y(_02828_)
  );
  sg13g2_o21ai_1 _13047_ (
    .A1(_02819_),
    .A2(_02828_),
    .B1(_00114_),
    .Y(_02829_)
  );
  sg13g2_a21oi_1 _13048_ (
    .A1(_01587_),
    .A2(_02107_),
    .B1(_01192_),
    .Y(_02830_)
  );
  sg13g2_nor2_1 _13049_ (
    .A(addr_i_4_),
    .B(_02830_),
    .Y(_02831_)
  );
  sg13g2_a21oi_1 _13050_ (
    .A1(addr_i_3_),
    .A2(_04384_),
    .B1(_05280_),
    .Y(_02833_)
  );
  sg13g2_o21ai_1 _13051_ (
    .A1(_02297_),
    .A2(_02833_),
    .B1(_02437_),
    .Y(_02834_)
  );
  sg13g2_a21o_1 _13052_ (
    .A1(_01738_),
    .A2(_07072_),
    .B1(addr_i_3_),
    .X(_02835_)
  );
  sg13g2_a21oi_1 _13053_ (
    .A1(_01462_),
    .A2(_02835_),
    .B1(addr_i_5_),
    .Y(_02836_)
  );
  sg13g2_or3_1 _13054_ (
    .A(_02831_),
    .B(_02834_),
    .C(_02836_),
    .X(_02837_)
  );
  sg13g2_nand2_1 _13055_ (
    .A(_01652_),
    .B(_00770_),
    .Y(_02838_)
  );
  sg13g2_a21oi_1 _13056_ (
    .A1(_00375_),
    .A2(_05258_),
    .B1(_02294_),
    .Y(_02839_)
  );
  sg13g2_nand2_1 _13057_ (
    .A(addr_i_3_),
    .B(_05689_),
    .Y(_02840_)
  );
  sg13g2_a21oi_1 _13058_ (
    .A1(_02304_),
    .A2(_02840_),
    .B1(_00899_),
    .Y(_02841_)
  );
  sg13g2_a22oi_1 _13059_ (
    .A1(_02838_),
    .A2(_02839_),
    .B1(_02841_),
    .B2(_00367_),
    .Y(_02842_)
  );
  sg13g2_a21oi_1 _13060_ (
    .A1(_02837_),
    .A2(_02842_),
    .B1(_06652_),
    .Y(_02844_)
  );
  sg13g2_nand2_1 _13061_ (
    .A(_02829_),
    .B(_02844_),
    .Y(_02845_)
  );
  sg13g2_nand4_1 _13062_ (
    .A(addr_i_11_),
    .B(_02767_),
    .C(_02814_),
    .D(_02845_),
    .Y(_02846_)
  );
  sg13g2_a21oi_1 _13063_ (
    .A1(_00245_),
    .A2(_00714_),
    .B1(_05269_),
    .Y(_02847_)
  );
  sg13g2_nor2_1 _13064_ (
    .A(addr_i_3_),
    .B(_00679_),
    .Y(_02848_)
  );
  sg13g2_o21ai_1 _13065_ (
    .A1(_02847_),
    .A2(_02848_),
    .B1(addr_i_4_),
    .Y(_02849_)
  );
  sg13g2_nor2_1 _13066_ (
    .A(addr_i_4_),
    .B(_04086_),
    .Y(_02850_)
  );
  sg13g2_a21oi_1 _13067_ (
    .A1(addr_i_4_),
    .A2(_00441_),
    .B1(addr_i_3_),
    .Y(_02851_)
  );
  sg13g2_o21ai_1 _13068_ (
    .A1(_02850_),
    .A2(_02851_),
    .B1(addr_i_7_),
    .Y(_02852_)
  );
  sg13g2_nand3_1 _13069_ (
    .A(_08022_),
    .B(_02849_),
    .C(_02852_),
    .Y(_02853_)
  );
  sg13g2_nand2_1 _13070_ (
    .A(addr_i_6_),
    .B(_02853_),
    .Y(_02855_)
  );
  sg13g2_o21ai_1 _13071_ (
    .A1(_00401_),
    .A2(_02494_),
    .B1(_09474_),
    .Y(_02856_)
  );
  sg13g2_a21oi_1 _13072_ (
    .A1(_02855_),
    .A2(_02856_),
    .B1(addr_i_8_),
    .Y(_02857_)
  );
  sg13g2_nand2_1 _13073_ (
    .A(addr_i_2_),
    .B(_06077_),
    .Y(_02858_)
  );
  sg13g2_o21ai_1 _13074_ (
    .A1(addr_i_4_),
    .A2(_02858_),
    .B1(_00353_),
    .Y(_02859_)
  );
  sg13g2_nand3_1 _13075_ (
    .A(addr_i_3_),
    .B(_01354_),
    .C(_02187_),
    .Y(_02860_)
  );
  sg13g2_o21ai_1 _13076_ (
    .A1(addr_i_3_),
    .A2(_02859_),
    .B1(_02860_),
    .Y(_02861_)
  );
  sg13g2_a22oi_1 _13077_ (
    .A1(_09483_),
    .A2(_01376_),
    .B1(_04672_),
    .B2(_01746_),
    .Y(_02862_)
  );
  sg13g2_nand4_1 _13078_ (
    .A(addr_i_6_),
    .B(_09105_),
    .C(_01118_),
    .D(_01287_),
    .Y(_02863_)
  );
  sg13g2_nand2_1 _13079_ (
    .A(_04119_),
    .B(_00008_),
    .Y(_02864_)
  );
  sg13g2_nand4_1 _13080_ (
    .A(_06717_),
    .B(_01118_),
    .C(_00872_),
    .D(_02864_),
    .Y(_02866_)
  );
  sg13g2_nand3_1 _13081_ (
    .A(addr_i_9_),
    .B(_02863_),
    .C(_02866_),
    .Y(_02867_)
  );
  sg13g2_a22oi_1 _13082_ (
    .A1(_01861_),
    .A2(_02861_),
    .B1(_02862_),
    .B2(_02867_),
    .Y(_02868_)
  );
  sg13g2_nor2b_1 _13083_ (
    .A(_02857_),
    .B_N(_02868_),
    .Y(_02869_)
  );
  sg13g2_a21oi_1 _13084_ (
    .A1(_02271_),
    .A2(_00591_),
    .B1(_07425_),
    .Y(_02870_)
  );
  sg13g2_nand2_1 _13085_ (
    .A(_08056_),
    .B(_02289_),
    .Y(_02871_)
  );
  sg13g2_o21ai_1 _13086_ (
    .A1(addr_i_4_),
    .A2(_02870_),
    .B1(_02871_),
    .Y(_02872_)
  );
  sg13g2_nor2_1 _13087_ (
    .A(_00547_),
    .B(_01197_),
    .Y(_02873_)
  );
  sg13g2_nand2_1 _13088_ (
    .A(addr_i_5_),
    .B(_07160_),
    .Y(_02874_)
  );
  sg13g2_a21oi_1 _13089_ (
    .A1(_01791_),
    .A2(_02874_),
    .B1(addr_i_3_),
    .Y(_02875_)
  );
  sg13g2_o21ai_1 _13090_ (
    .A1(_02873_),
    .A2(_02875_),
    .B1(_03930_),
    .Y(_02877_)
  );
  sg13g2_a21oi_1 _13091_ (
    .A1(_00007_),
    .A2(_02089_),
    .B1(_02076_),
    .Y(_02878_)
  );
  sg13g2_nor2_1 _13092_ (
    .A(addr_i_4_),
    .B(_02878_),
    .Y(_02879_)
  );
  sg13g2_nand2_1 _13093_ (
    .A(addr_i_7_),
    .B(_02076_),
    .Y(_02880_)
  );
  sg13g2_o21ai_1 _13094_ (
    .A1(_00454_),
    .A2(_08100_),
    .B1(addr_i_3_),
    .Y(_02881_)
  );
  sg13g2_a21oi_1 _13095_ (
    .A1(_04296_),
    .A2(_02881_),
    .B1(_04251_),
    .Y(_02882_)
  );
  sg13g2_a22oi_1 _13096_ (
    .A1(_07547_),
    .A2(_02880_),
    .B1(_02882_),
    .B2(_08399_),
    .Y(_02883_)
  );
  sg13g2_a22oi_1 _13097_ (
    .A1(_02877_),
    .A2(_02879_),
    .B1(_00367_),
    .B2(_02883_),
    .Y(_02884_)
  );
  sg13g2_a21oi_1 _13098_ (
    .A1(_00277_),
    .A2(_02872_),
    .B1(_02884_),
    .Y(_02885_)
  );
  sg13g2_o21ai_1 _13099_ (
    .A1(addr_i_9_),
    .A2(_02885_),
    .B1(_00511_),
    .Y(_02886_)
  );
  sg13g2_nand2_1 _13100_ (
    .A(_01208_),
    .B(_09478_),
    .Y(_02888_)
  );
  sg13g2_a22oi_1 _13101_ (
    .A1(_02796_),
    .A2(_02888_),
    .B1(_00192_),
    .B2(_05822_),
    .Y(_02889_)
  );
  sg13g2_nand2_1 _13102_ (
    .A(_02799_),
    .B(_01636_),
    .Y(_02890_)
  );
  sg13g2_nor2_1 _13103_ (
    .A(_03743_),
    .B(_00008_),
    .Y(_02891_)
  );
  sg13g2_a22oi_1 _13104_ (
    .A1(_01450_),
    .A2(_02890_),
    .B1(_02891_),
    .B2(addr_i_7_),
    .Y(_02892_)
  );
  sg13g2_nor2_1 _13105_ (
    .A(_02889_),
    .B(_02892_),
    .Y(_02893_)
  );
  sg13g2_nand2_1 _13106_ (
    .A(_08266_),
    .B(_01234_),
    .Y(_02894_)
  );
  sg13g2_nand2_1 _13107_ (
    .A(_00915_),
    .B(_08111_),
    .Y(_02895_)
  );
  sg13g2_a21oi_1 _13108_ (
    .A1(_01786_),
    .A2(_02895_),
    .B1(addr_i_7_),
    .Y(_02896_)
  );
  sg13g2_a22oi_1 _13109_ (
    .A1(_02277_),
    .A2(_02894_),
    .B1(_02896_),
    .B2(_00029_),
    .Y(_02897_)
  );
  sg13g2_o21ai_1 _13110_ (
    .A1(addr_i_2_),
    .A2(_02897_),
    .B1(addr_i_8_),
    .Y(_02899_)
  );
  sg13g2_nand4_1 _13111_ (
    .A(addr_i_4_),
    .B(_06895_),
    .C(_00315_),
    .D(_01514_),
    .Y(_02900_)
  );
  sg13g2_a21oi_1 _13112_ (
    .A1(_07790_),
    .A2(_00943_),
    .B1(addr_i_4_),
    .Y(_02901_)
  );
  sg13g2_a22oi_1 _13113_ (
    .A1(_07824_),
    .A2(_00561_),
    .B1(_00860_),
    .B2(_02901_),
    .Y(_02902_)
  );
  sg13g2_a21oi_1 _13114_ (
    .A1(_09478_),
    .A2(_00872_),
    .B1(addr_i_6_),
    .Y(_02903_)
  );
  sg13g2_nor2_1 _13115_ (
    .A(_08830_),
    .B(_02903_),
    .Y(_02904_)
  );
  sg13g2_a21oi_1 _13116_ (
    .A1(_02900_),
    .A2(_02902_),
    .B1(_02904_),
    .Y(_02905_)
  );
  sg13g2_o21ai_1 _13117_ (
    .A1(_02893_),
    .A2(_02899_),
    .B1(_02905_),
    .Y(_02906_)
  );
  sg13g2_nor3_1 _13118_ (
    .A(addr_i_2_),
    .B(_01473_),
    .C(_01519_),
    .Y(_02907_)
  );
  sg13g2_o21ai_1 _13119_ (
    .A1(_01002_),
    .A2(_02907_),
    .B1(addr_i_7_),
    .Y(_02908_)
  );
  sg13g2_o21ai_1 _13120_ (
    .A1(_06563_),
    .A2(_02652_),
    .B1(_00293_),
    .Y(_02910_)
  );
  sg13g2_a21oi_1 _13121_ (
    .A1(_01410_),
    .A2(_02910_),
    .B1(addr_i_4_),
    .Y(_02911_)
  );
  sg13g2_a22oi_1 _13122_ (
    .A1(_00301_),
    .A2(_00031_),
    .B1(_02911_),
    .B2(_00629_),
    .Y(_02912_)
  );
  sg13g2_o21ai_1 _13123_ (
    .A1(_07337_),
    .A2(_00258_),
    .B1(_07625_),
    .Y(_02913_)
  );
  sg13g2_a21oi_1 _13124_ (
    .A1(addr_i_6_),
    .A2(_02913_),
    .B1(_07614_),
    .Y(_02914_)
  );
  sg13g2_a22oi_1 _13125_ (
    .A1(_01240_),
    .A2(_02567_),
    .B1(_01819_),
    .B2(_00802_),
    .Y(_02915_)
  );
  sg13g2_a22oi_1 _13126_ (
    .A1(_02908_),
    .A2(_02912_),
    .B1(_02914_),
    .B2(_02915_),
    .Y(_02916_)
  );
  sg13g2_nor2_1 _13127_ (
    .A(_02221_),
    .B(_02916_),
    .Y(_02917_)
  );
  sg13g2_a22oi_1 _13128_ (
    .A1(_01176_),
    .A2(_02906_),
    .B1(_02917_),
    .B2(addr_i_11_),
    .Y(_02918_)
  );
  sg13g2_o21ai_1 _13129_ (
    .A1(_02869_),
    .A2(_02886_),
    .B1(_02918_),
    .Y(_02919_)
  );
  sg13g2_nand3_1 _13130_ (
    .A(_02251_),
    .B(_02846_),
    .C(_02919_),
    .Y(_02921_)
  );
  sg13g2_o21ai_1 _13131_ (
    .A1(_02716_),
    .A2(_02741_),
    .B1(_02921_),
    .Y(data_o_16_)
  );
  sg13g2_a21oi_1 _13132_ (
    .A1(_00104_),
    .A2(_00228_),
    .B1(_00479_),
    .Y(_02922_)
  );
  sg13g2_a21oi_1 _13133_ (
    .A1(_05457_),
    .A2(_01084_),
    .B1(addr_i_3_),
    .Y(_02923_)
  );
  sg13g2_nor3_1 _13134_ (
    .A(_00548_),
    .B(_02922_),
    .C(_02923_),
    .Y(_02924_)
  );
  sg13g2_nor2_1 _13135_ (
    .A(addr_i_3_),
    .B(_01375_),
    .Y(_02925_)
  );
  sg13g2_o21ai_1 _13136_ (
    .A1(_01456_),
    .A2(_02925_),
    .B1(_09138_),
    .Y(_02926_)
  );
  sg13g2_nand3b_1 _13137_ (
    .A_N(_02924_),
    .B(addr_i_8_),
    .C(_02926_),
    .Y(_02927_)
  );
  sg13g2_nand2_1 _13138_ (
    .A(_00462_),
    .B(_05678_),
    .Y(_02928_)
  );
  sg13g2_a22oi_1 _13139_ (
    .A1(addr_i_3_),
    .A2(_02928_),
    .B1(_01660_),
    .B2(_00007_),
    .Y(_02929_)
  );
  sg13g2_nand2_1 _13140_ (
    .A(addr_i_3_),
    .B(_02472_),
    .Y(_02931_)
  );
  sg13g2_a21oi_1 _13141_ (
    .A1(_01897_),
    .A2(_02931_),
    .B1(_00548_),
    .Y(_02932_)
  );
  sg13g2_or3_1 _13142_ (
    .A(addr_i_8_),
    .B(_02929_),
    .C(_02932_),
    .X(_02933_)
  );
  sg13g2_nand2_1 _13143_ (
    .A(_02927_),
    .B(_02933_),
    .Y(_02934_)
  );
  sg13g2_nor2_1 _13144_ (
    .A(addr_i_3_),
    .B(_00725_),
    .Y(_02935_)
  );
  sg13g2_o21ai_1 _13145_ (
    .A1(_01500_),
    .A2(_02935_),
    .B1(addr_i_4_),
    .Y(_02936_)
  );
  sg13g2_a21oi_1 _13146_ (
    .A1(_06884_),
    .A2(_01588_),
    .B1(_05856_),
    .Y(_02937_)
  );
  sg13g2_o21ai_1 _13147_ (
    .A1(_01493_),
    .A2(_02937_),
    .B1(addr_i_2_),
    .Y(_02938_)
  );
  sg13g2_nand3_1 _13148_ (
    .A(_01182_),
    .B(_02936_),
    .C(_02938_),
    .Y(_02939_)
  );
  sg13g2_o21ai_1 _13149_ (
    .A1(_02933_),
    .A2(_02939_),
    .B1(_05203_),
    .Y(_02940_)
  );
  sg13g2_nor2_1 _13150_ (
    .A(addr_i_3_),
    .B(_06541_),
    .Y(_02942_)
  );
  sg13g2_a21oi_1 _13151_ (
    .A1(addr_i_4_),
    .A2(_04075_),
    .B1(_04086_),
    .Y(_02943_)
  );
  sg13g2_nand2_1 _13152_ (
    .A(addr_i_6_),
    .B(_02304_),
    .Y(_02944_)
  );
  sg13g2_o21ai_1 _13153_ (
    .A1(addr_i_6_),
    .A2(_02943_),
    .B1(_02944_),
    .Y(_02945_)
  );
  sg13g2_a221oi_1 _13154_ (
    .A1(_09483_),
    .A2(_02942_),
    .B1(_02945_),
    .B2(addr_i_3_),
    .C1(_02927_),
    .Y(_02946_)
  );
  sg13g2_a22oi_1 _13155_ (
    .A1(addr_i_7_),
    .A2(_02934_),
    .B1(_02940_),
    .B2(_02946_),
    .Y(_02947_)
  );
  sg13g2_nand2_1 _13156_ (
    .A(_00581_),
    .B(_06851_),
    .Y(_02948_)
  );
  sg13g2_nor2_1 _13157_ (
    .A(_00534_),
    .B(_06032_),
    .Y(_02949_)
  );
  sg13g2_a22oi_1 _13158_ (
    .A1(_00626_),
    .A2(_02948_),
    .B1(_02949_),
    .B2(_08487_),
    .Y(_02950_)
  );
  sg13g2_o21ai_1 _13159_ (
    .A1(_03150_),
    .A2(_00416_),
    .B1(addr_i_3_),
    .Y(_02951_)
  );
  sg13g2_nand2_1 _13160_ (
    .A(addr_i_4_),
    .B(_09382_),
    .Y(_02953_)
  );
  sg13g2_nor2_1 _13161_ (
    .A(addr_i_3_),
    .B(_05966_),
    .Y(_02954_)
  );
  sg13g2_nand3_1 _13162_ (
    .A(_01050_),
    .B(_02953_),
    .C(_02954_),
    .Y(_02955_)
  );
  sg13g2_nand3_1 _13163_ (
    .A(_05302_),
    .B(addr_i_6_),
    .C(_02755_),
    .Y(_02956_)
  );
  sg13g2_nand3_1 _13164_ (
    .A(addr_i_3_),
    .B(_02052_),
    .C(_02956_),
    .Y(_02957_)
  );
  sg13g2_a21oi_1 _13165_ (
    .A1(_02955_),
    .A2(_02957_),
    .B1(_01082_),
    .Y(_02958_)
  );
  sg13g2_or2_1 _13166_ (
    .A(_07348_),
    .B(_01777_),
    .X(_02959_)
  );
  sg13g2_a221oi_1 _13167_ (
    .A1(_00073_),
    .A2(_00136_),
    .B1(_02959_),
    .B2(_01282_),
    .C1(_01391_),
    .Y(_02960_)
  );
  sg13g2_a22oi_1 _13168_ (
    .A1(_02950_),
    .A2(_02951_),
    .B1(_02958_),
    .B2(_02960_),
    .Y(_02961_)
  );
  sg13g2_nand2_1 _13169_ (
    .A(addr_i_3_),
    .B(_00666_),
    .Y(_02962_)
  );
  sg13g2_a21oi_1 _13170_ (
    .A1(_00595_),
    .A2(_02962_),
    .B1(addr_i_2_),
    .Y(_02964_)
  );
  sg13g2_nand2_1 _13171_ (
    .A(addr_i_4_),
    .B(_05435_),
    .Y(_02965_)
  );
  sg13g2_nand3_1 _13172_ (
    .A(_00084_),
    .B(_07790_),
    .C(_00211_),
    .Y(_02966_)
  );
  sg13g2_o21ai_1 _13173_ (
    .A1(_02964_),
    .A2(_02965_),
    .B1(_02966_),
    .Y(_02967_)
  );
  sg13g2_nand2_1 _13174_ (
    .A(_00277_),
    .B(_02967_),
    .Y(_02968_)
  );
  sg13g2_a21oi_1 _13175_ (
    .A1(_02961_),
    .A2(_02968_),
    .B1(_01211_),
    .Y(_02969_)
  );
  sg13g2_o21ai_1 _13176_ (
    .A1(_08100_),
    .A2(_07105_),
    .B1(addr_i_4_),
    .Y(_02970_)
  );
  sg13g2_nand3_1 _13177_ (
    .A(addr_i_3_),
    .B(_02661_),
    .C(_02970_),
    .Y(_02971_)
  );
  sg13g2_o21ai_1 _13178_ (
    .A1(addr_i_7_),
    .A2(_07636_),
    .B1(_01113_),
    .Y(_02972_)
  );
  sg13g2_nand2_1 _13179_ (
    .A(_07668_),
    .B(_02972_),
    .Y(_02973_)
  );
  sg13g2_a21oi_1 _13180_ (
    .A1(_02971_),
    .A2(_02973_),
    .B1(_08708_),
    .Y(_02975_)
  );
  sg13g2_buf_1 _13181_ (
    .A(_00086_),
    .X(_02976_)
  );
  sg13g2_a21oi_1 _13182_ (
    .A1(_01592_),
    .A2(_08221_),
    .B1(_01120_),
    .Y(_02977_)
  );
  sg13g2_a22oi_1 _13183_ (
    .A1(_02976_),
    .A2(_07503_),
    .B1(_02977_),
    .B2(addr_i_5_),
    .Y(_02978_)
  );
  sg13g2_or2_1 _13184_ (
    .A(_02975_),
    .B(_02978_),
    .X(_02979_)
  );
  sg13g2_nor2_1 _13185_ (
    .A(addr_i_5_),
    .B(_00099_),
    .Y(_02980_)
  );
  sg13g2_o21ai_1 _13186_ (
    .A1(_05025_),
    .A2(_02980_),
    .B1(addr_i_6_),
    .Y(_02981_)
  );
  sg13g2_a21oi_1 _13187_ (
    .A1(_04296_),
    .A2(_02981_),
    .B1(_00565_),
    .Y(_02982_)
  );
  sg13g2_nor2_1 _13188_ (
    .A(_02196_),
    .B(_02558_),
    .Y(_02983_)
  );
  sg13g2_nor4_1 _13189_ (
    .A(addr_i_8_),
    .B(_04506_),
    .C(_02982_),
    .D(_02983_),
    .Y(_02984_)
  );
  sg13g2_a21oi_1 _13190_ (
    .A1(_00870_),
    .A2(_01708_),
    .B1(addr_i_7_),
    .Y(_02986_)
  );
  sg13g2_nand2_1 _13191_ (
    .A(_00454_),
    .B(_07492_),
    .Y(_02987_)
  );
  sg13g2_a21oi_1 _13192_ (
    .A1(_01543_),
    .A2(_02987_),
    .B1(addr_i_6_),
    .Y(_02988_)
  );
  sg13g2_nor3_1 _13193_ (
    .A(_01577_),
    .B(_02986_),
    .C(_02988_),
    .Y(_02989_)
  );
  sg13g2_buf_1 _13194_ (
    .A(_08156_),
    .X(_02990_)
  );
  sg13g2_nor3_1 _13195_ (
    .A(_02990_),
    .B(addr_i_6_),
    .C(_00001_),
    .Y(_02991_)
  );
  sg13g2_a21oi_1 _13196_ (
    .A1(_01527_),
    .A2(_01886_),
    .B1(addr_i_7_),
    .Y(_02992_)
  );
  sg13g2_o21ai_1 _13197_ (
    .A1(_02991_),
    .A2(_02992_),
    .B1(addr_i_4_),
    .Y(_02993_)
  );
  sg13g2_nand2_1 _13198_ (
    .A(_00342_),
    .B(_00624_),
    .Y(_02994_)
  );
  sg13g2_o21ai_1 _13199_ (
    .A1(_00384_),
    .A2(_02490_),
    .B1(_03919_),
    .Y(_02995_)
  );
  sg13g2_a21o_1 _13200_ (
    .A1(_02994_),
    .A2(_02995_),
    .B1(_04251_),
    .X(_02997_)
  );
  sg13g2_nand3_1 _13201_ (
    .A(_02989_),
    .B(_02993_),
    .C(_02997_),
    .Y(_02998_)
  );
  sg13g2_a221oi_1 _13202_ (
    .A1(_02979_),
    .A2(_02984_),
    .B1(_02998_),
    .B2(addr_i_8_),
    .C1(addr_i_9_),
    .Y(_02999_)
  );
  sg13g2_inv_1 _13203_ (
    .A(_02999_),
    .Y(_03000_)
  );
  sg13g2_nor3_1 _13204_ (
    .A(addr_i_2_),
    .B(_00001_),
    .C(_05645_),
    .Y(_03001_)
  );
  sg13g2_nand3_1 _13205_ (
    .A(_08410_),
    .B(_02994_),
    .C(_00250_),
    .Y(_03002_)
  );
  sg13g2_nor2b_1 _13206_ (
    .A(_03001_),
    .B_N(_03002_),
    .Y(_03003_)
  );
  sg13g2_nor2_1 _13207_ (
    .A(_05722_),
    .B(_06530_),
    .Y(_03004_)
  );
  sg13g2_nor3_1 _13208_ (
    .A(addr_i_4_),
    .B(_00990_),
    .C(_02976_),
    .Y(_03005_)
  );
  sg13g2_a22oi_1 _13209_ (
    .A1(addr_i_4_),
    .A2(_03004_),
    .B1(_03005_),
    .B2(addr_i_3_),
    .Y(_03006_)
  );
  sg13g2_o21ai_1 _13210_ (
    .A1(_07348_),
    .A2(_09502_),
    .B1(_01308_),
    .Y(_03008_)
  );
  sg13g2_nand2_1 _13211_ (
    .A(_00324_),
    .B(_03008_),
    .Y(_03009_)
  );
  sg13g2_a22oi_1 _13212_ (
    .A1(addr_i_3_),
    .A2(_03003_),
    .B1(_03006_),
    .B2(_03009_),
    .Y(_03010_)
  );
  sg13g2_nand2b_1 _13213_ (
    .A_N(_03010_),
    .B(_00469_),
    .Y(_03011_)
  );
  sg13g2_nor2_1 _13214_ (
    .A(_07049_),
    .B(_00923_),
    .Y(_03012_)
  );
  sg13g2_o21ai_1 _13215_ (
    .A1(_00605_),
    .A2(_03012_),
    .B1(_01120_),
    .Y(_03013_)
  );
  sg13g2_o21ai_1 _13216_ (
    .A1(addr_i_3_),
    .A2(_02342_),
    .B1(_03013_),
    .Y(_03014_)
  );
  sg13g2_o21ai_1 _13217_ (
    .A1(_00700_),
    .A2(_09448_),
    .B1(_01290_),
    .Y(_03015_)
  );
  sg13g2_a221oi_1 _13218_ (
    .A1(addr_i_2_),
    .A2(_03014_),
    .B1(_03015_),
    .B2(addr_i_4_),
    .C1(addr_i_7_),
    .Y(_03016_)
  );
  sg13g2_o21ai_1 _13219_ (
    .A1(_00840_),
    .A2(_00503_),
    .B1(_01528_),
    .Y(_03017_)
  );
  sg13g2_o21ai_1 _13220_ (
    .A1(_01459_),
    .A2(_00861_),
    .B1(addr_i_4_),
    .Y(_03019_)
  );
  sg13g2_a21oi_1 _13221_ (
    .A1(_03017_),
    .A2(_03019_),
    .B1(_02759_),
    .Y(_03020_)
  );
  sg13g2_xnor2_1 _13222_ (
    .A(addr_i_5_),
    .B(_00711_),
    .Y(_03021_)
  );
  sg13g2_nand2_1 _13223_ (
    .A(_09497_),
    .B(_00712_),
    .Y(_03022_)
  );
  sg13g2_o21ai_1 _13224_ (
    .A1(addr_i_4_),
    .A2(_03021_),
    .B1(_03022_),
    .Y(_03023_)
  );
  sg13g2_o21ai_1 _13225_ (
    .A1(_00548_),
    .A2(_03023_),
    .B1(addr_i_8_),
    .Y(_03024_)
  );
  sg13g2_or3_1 _13226_ (
    .A(_03016_),
    .B(_03020_),
    .C(_03024_),
    .X(_03025_)
  );
  sg13g2_nand3_1 _13227_ (
    .A(addr_i_9_),
    .B(_03011_),
    .C(_03025_),
    .Y(_03026_)
  );
  sg13g2_a21oi_1 _13228_ (
    .A1(_03000_),
    .A2(_03026_),
    .B1(addr_i_10_),
    .Y(_03027_)
  );
  sg13g2_nor4_1 _13229_ (
    .A(addr_i_11_),
    .B(_02947_),
    .C(_02969_),
    .D(_03027_),
    .Y(_03028_)
  );
  sg13g2_nor2_1 _13230_ (
    .A(addr_i_4_),
    .B(_00588_),
    .Y(_03030_)
  );
  sg13g2_a21oi_1 _13231_ (
    .A1(_03238_),
    .A2(_01656_),
    .B1(_03030_),
    .Y(_03031_)
  );
  sg13g2_nor3_1 _13232_ (
    .A(addr_i_3_),
    .B(addr_i_4_),
    .C(addr_i_5_),
    .Y(_03032_)
  );
  sg13g2_buf_1 _13233_ (
    .A(_03032_),
    .X(_03033_)
  );
  sg13g2_o21ai_1 _13234_ (
    .A1(_03033_),
    .A2(_00266_),
    .B1(addr_i_6_),
    .Y(_03034_)
  );
  sg13g2_o21ai_1 _13235_ (
    .A1(addr_i_3_),
    .A2(_01282_),
    .B1(_02694_),
    .Y(_03035_)
  );
  sg13g2_a21oi_1 _13236_ (
    .A1(_01815_),
    .A2(_01514_),
    .B1(addr_i_2_),
    .Y(_03036_)
  );
  sg13g2_a22oi_1 _13237_ (
    .A1(addr_i_4_),
    .A2(_03035_),
    .B1(_03036_),
    .B2(addr_i_7_),
    .Y(_03037_)
  );
  sg13g2_a221oi_1 _13238_ (
    .A1(addr_i_7_),
    .A2(_01656_),
    .B1(_03034_),
    .B2(_03037_),
    .C1(_01612_),
    .Y(_03038_)
  );
  sg13g2_nor2_1 _13239_ (
    .A(_02371_),
    .B(_02459_),
    .Y(_03039_)
  );
  sg13g2_a21oi_1 _13240_ (
    .A1(_03424_),
    .A2(_00391_),
    .B1(addr_i_3_),
    .Y(_03041_)
  );
  sg13g2_o21ai_1 _13241_ (
    .A1(_03039_),
    .A2(_03041_),
    .B1(_00388_),
    .Y(_03042_)
  );
  sg13g2_a21oi_1 _13242_ (
    .A1(_00007_),
    .A2(_02577_),
    .B1(_02744_),
    .Y(_03043_)
  );
  sg13g2_o21ai_1 _13243_ (
    .A1(addr_i_2_),
    .A2(_02091_),
    .B1(_03043_),
    .Y(_03044_)
  );
  sg13g2_nor2_1 _13244_ (
    .A(addr_i_6_),
    .B(_08885_),
    .Y(_03045_)
  );
  sg13g2_nand2_1 _13245_ (
    .A(_00463_),
    .B(_06884_),
    .Y(_03046_)
  );
  sg13g2_o21ai_1 _13246_ (
    .A1(_02387_),
    .A2(_03045_),
    .B1(_03046_),
    .Y(_03047_)
  );
  sg13g2_nand3_1 _13247_ (
    .A(addr_i_7_),
    .B(_00138_),
    .C(_00287_),
    .Y(_03048_)
  );
  sg13g2_o21ai_1 _13248_ (
    .A1(addr_i_7_),
    .A2(_03047_),
    .B1(_03048_),
    .Y(_03049_)
  );
  sg13g2_nand2_1 _13249_ (
    .A(addr_i_4_),
    .B(_03049_),
    .Y(_03050_)
  );
  sg13g2_and4_1 _13250_ (
    .A(_00423_),
    .B(_03042_),
    .C(_03044_),
    .D(_03050_),
    .X(_03052_)
  );
  sg13g2_a22oi_1 _13251_ (
    .A1(addr_i_9_),
    .A2(_03031_),
    .B1(_03038_),
    .B2(_03052_),
    .Y(_03053_)
  );
  sg13g2_o21ai_1 _13252_ (
    .A1(_02744_),
    .A2(_09260_),
    .B1(_02136_),
    .Y(_03054_)
  );
  sg13g2_a21oi_1 _13253_ (
    .A1(_01350_),
    .A2(_03054_),
    .B1(_01640_),
    .Y(_03055_)
  );
  sg13g2_o21ai_1 _13254_ (
    .A1(addr_i_10_),
    .A2(_03053_),
    .B1(_03055_),
    .Y(_03056_)
  );
  sg13g2_nand2_1 _13255_ (
    .A(addr_i_12_),
    .B(_03056_),
    .Y(_03057_)
  );
  sg13g2_nand2_1 _13256_ (
    .A(_02089_),
    .B(_01618_),
    .Y(_03058_)
  );
  sg13g2_nor2_1 _13257_ (
    .A(_00695_),
    .B(_01128_),
    .Y(_03059_)
  );
  sg13g2_a22oi_1 _13258_ (
    .A1(addr_i_4_),
    .A2(_03058_),
    .B1(_03059_),
    .B2(_02530_),
    .Y(_03060_)
  );
  sg13g2_a21oi_1 _13259_ (
    .A1(addr_i_4_),
    .A2(_01066_),
    .B1(_07636_),
    .Y(_03061_)
  );
  sg13g2_a221oi_1 _13260_ (
    .A1(_00818_),
    .A2(_01421_),
    .B1(_03061_),
    .B2(_00377_),
    .C1(addr_i_3_),
    .Y(_03063_)
  );
  sg13g2_a21oi_1 _13261_ (
    .A1(_00500_),
    .A2(_05645_),
    .B1(addr_i_8_),
    .Y(_03064_)
  );
  sg13g2_o21ai_1 _13262_ (
    .A1(_03060_),
    .A2(_03063_),
    .B1(_03064_),
    .Y(_03065_)
  );
  sg13g2_nor2_1 _13263_ (
    .A(_01301_),
    .B(_00254_),
    .Y(_03066_)
  );
  sg13g2_a21oi_1 _13264_ (
    .A1(addr_i_4_),
    .A2(_00138_),
    .B1(_00778_),
    .Y(_03067_)
  );
  sg13g2_o21ai_1 _13265_ (
    .A1(_03066_),
    .A2(_03067_),
    .B1(addr_i_3_),
    .Y(_03068_)
  );
  sg13g2_o21ai_1 _13266_ (
    .A1(_00959_),
    .A2(_00503_),
    .B1(_02118_),
    .Y(_03069_)
  );
  sg13g2_nor2_1 _13267_ (
    .A(addr_i_4_),
    .B(_05756_),
    .Y(_03070_)
  );
  sg13g2_nand2_1 _13268_ (
    .A(_01970_),
    .B(_03070_),
    .Y(_03071_)
  );
  sg13g2_o21ai_1 _13269_ (
    .A1(_02330_),
    .A2(_02361_),
    .B1(addr_i_4_),
    .Y(_03072_)
  );
  sg13g2_a21o_1 _13270_ (
    .A1(_03071_),
    .A2(_03072_),
    .B1(addr_i_7_),
    .X(_03074_)
  );
  sg13g2_nand4_1 _13271_ (
    .A(addr_i_8_),
    .B(_03068_),
    .C(_03069_),
    .D(_03074_),
    .Y(_03075_)
  );
  sg13g2_nand3_1 _13272_ (
    .A(addr_i_9_),
    .B(_03065_),
    .C(_03075_),
    .Y(_03076_)
  );
  sg13g2_nor2_1 _13273_ (
    .A(_06298_),
    .B(_07270_),
    .Y(_03077_)
  );
  sg13g2_o21ai_1 _13274_ (
    .A1(addr_i_4_),
    .A2(_03077_),
    .B1(_09039_),
    .Y(_03078_)
  );
  sg13g2_o21ai_1 _13275_ (
    .A1(_01954_),
    .A2(_00346_),
    .B1(addr_i_2_),
    .Y(_03079_)
  );
  sg13g2_nand3_1 _13276_ (
    .A(addr_i_6_),
    .B(_01473_),
    .C(_03079_),
    .Y(_03080_)
  );
  sg13g2_o21ai_1 _13277_ (
    .A1(addr_i_6_),
    .A2(_03078_),
    .B1(_03080_),
    .Y(_03081_)
  );
  sg13g2_o21ai_1 _13278_ (
    .A1(_01024_),
    .A2(_09215_),
    .B1(addr_i_3_),
    .Y(_03082_)
  );
  sg13g2_a21oi_1 _13279_ (
    .A1(addr_i_6_),
    .A2(_00692_),
    .B1(_01473_),
    .Y(_03083_)
  );
  sg13g2_nand2_1 _13280_ (
    .A(_06862_),
    .B(_02462_),
    .Y(_03085_)
  );
  sg13g2_nand3_1 _13281_ (
    .A(_00339_),
    .B(_07934_),
    .C(_03085_),
    .Y(_03086_)
  );
  sg13g2_nor2_1 _13282_ (
    .A(_03083_),
    .B(_03086_),
    .Y(_03087_)
  );
  sg13g2_a221oi_1 _13283_ (
    .A1(_01666_),
    .A2(_03081_),
    .B1(_03082_),
    .B2(_03087_),
    .C1(addr_i_9_),
    .Y(_03088_)
  );
  sg13g2_nand2_1 _13284_ (
    .A(_00078_),
    .B(_05678_),
    .Y(_03089_)
  );
  sg13g2_a21o_1 _13285_ (
    .A1(addr_i_3_),
    .A2(_03089_),
    .B1(_01746_),
    .X(_03090_)
  );
  sg13g2_o21ai_1 _13286_ (
    .A1(_05258_),
    .A2(_01910_),
    .B1(addr_i_3_),
    .Y(_03091_)
  );
  sg13g2_a21oi_1 _13287_ (
    .A1(_08022_),
    .A2(_03091_),
    .B1(_00492_),
    .Y(_03092_)
  );
  sg13g2_a22oi_1 _13288_ (
    .A1(_01542_),
    .A2(_03090_),
    .B1(_03092_),
    .B2(addr_i_8_),
    .Y(_03093_)
  );
  sg13g2_o21ai_1 _13289_ (
    .A1(_02181_),
    .A2(_01659_),
    .B1(_00059_),
    .Y(_03094_)
  );
  sg13g2_a21oi_1 _13290_ (
    .A1(_00771_),
    .A2(_03094_),
    .B1(addr_i_6_),
    .Y(_03096_)
  );
  sg13g2_nor2_1 _13291_ (
    .A(_00080_),
    .B(_02583_),
    .Y(_03097_)
  );
  sg13g2_o21ai_1 _13292_ (
    .A1(_03096_),
    .A2(_03097_),
    .B1(addr_i_7_),
    .Y(_03098_)
  );
  sg13g2_nand2_1 _13293_ (
    .A(_03093_),
    .B(_03098_),
    .Y(_03099_)
  );
  sg13g2_a21oi_1 _13294_ (
    .A1(_03088_),
    .A2(_03099_),
    .B1(_01773_),
    .Y(_03100_)
  );
  sg13g2_a21oi_1 _13295_ (
    .A1(addr_i_2_),
    .A2(_01813_),
    .B1(_06099_),
    .Y(_03101_)
  );
  sg13g2_nor2_1 _13296_ (
    .A(_00726_),
    .B(_03101_),
    .Y(_03102_)
  );
  sg13g2_o21ai_1 _13297_ (
    .A1(_00278_),
    .A2(_09183_),
    .B1(addr_i_4_),
    .Y(_03103_)
  );
  sg13g2_o21ai_1 _13298_ (
    .A1(_01106_),
    .A2(_02376_),
    .B1(addr_i_6_),
    .Y(_03104_)
  );
  sg13g2_nand3_1 _13299_ (
    .A(addr_i_7_),
    .B(_03103_),
    .C(_03104_),
    .Y(_03105_)
  );
  sg13g2_o21ai_1 _13300_ (
    .A1(_03102_),
    .A2(_03105_),
    .B1(addr_i_8_),
    .Y(_03107_)
  );
  sg13g2_nand2_1 _13301_ (
    .A(_02020_),
    .B(_00252_),
    .Y(_03108_)
  );
  sg13g2_nand3_1 _13302_ (
    .A(addr_i_3_),
    .B(_00567_),
    .C(_03108_),
    .Y(_03109_)
  );
  sg13g2_buf_1 _13303_ (
    .A(_00835_),
    .X(_03110_)
  );
  sg13g2_nand3_1 _13304_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .C(_03110_),
    .Y(_03111_)
  );
  sg13g2_nor2_1 _13305_ (
    .A(_06386_),
    .B(_05335_),
    .Y(_03112_)
  );
  sg13g2_nand2_1 _13306_ (
    .A(_04108_),
    .B(_03112_),
    .Y(_03113_)
  );
  sg13g2_nand3_1 _13307_ (
    .A(_05867_),
    .B(_03111_),
    .C(_03113_),
    .Y(_03114_)
  );
  sg13g2_a21oi_1 _13308_ (
    .A1(_03109_),
    .A2(_03114_),
    .B1(addr_i_7_),
    .Y(_03115_)
  );
  sg13g2_nand2_1 _13309_ (
    .A(_04650_),
    .B(_02732_),
    .Y(_03116_)
  );
  sg13g2_o21ai_1 _13310_ (
    .A1(addr_i_6_),
    .A2(_00014_),
    .B1(addr_i_4_),
    .Y(_03118_)
  );
  sg13g2_a21oi_1 _13311_ (
    .A1(_00906_),
    .A2(_03118_),
    .B1(_02105_),
    .Y(_03119_)
  );
  sg13g2_a22oi_1 _13312_ (
    .A1(_00910_),
    .A2(_01264_),
    .B1(_03116_),
    .B2(_03119_),
    .Y(_03120_)
  );
  sg13g2_nor3_1 _13313_ (
    .A(addr_i_3_),
    .B(addr_i_5_),
    .C(_01014_),
    .Y(_03121_)
  );
  sg13g2_nor2_1 _13314_ (
    .A(_01112_),
    .B(_03121_),
    .Y(_03122_)
  );
  sg13g2_a21oi_1 _13315_ (
    .A1(_00736_),
    .A2(_00870_),
    .B1(addr_i_6_),
    .Y(_03123_)
  );
  sg13g2_a22oi_1 _13316_ (
    .A1(addr_i_3_),
    .A2(_01789_),
    .B1(_03123_),
    .B2(_08155_),
    .Y(_03124_)
  );
  sg13g2_a22oi_1 _13317_ (
    .A1(_00360_),
    .A2(_03122_),
    .B1(_03124_),
    .B2(_00860_),
    .Y(_03125_)
  );
  sg13g2_nor2_1 _13318_ (
    .A(_03120_),
    .B(_03125_),
    .Y(_03126_)
  );
  sg13g2_o21ai_1 _13319_ (
    .A1(_03107_),
    .A2(_03115_),
    .B1(_03126_),
    .Y(_03127_)
  );
  sg13g2_nand2_1 _13320_ (
    .A(_00914_),
    .B(_02799_),
    .Y(_03129_)
  );
  sg13g2_a21oi_1 _13321_ (
    .A1(addr_i_3_),
    .A2(_03129_),
    .B1(_01746_),
    .Y(_03130_)
  );
  sg13g2_nand2_1 _13322_ (
    .A(_05258_),
    .B(_07458_),
    .Y(_03131_)
  );
  sg13g2_nand2_1 _13323_ (
    .A(addr_i_6_),
    .B(_00713_),
    .Y(_03132_)
  );
  sg13g2_a21oi_1 _13324_ (
    .A1(_00581_),
    .A2(_00406_),
    .B1(_05856_),
    .Y(_03133_)
  );
  sg13g2_nor3_1 _13325_ (
    .A(_02261_),
    .B(_03132_),
    .C(_03133_),
    .Y(_03134_)
  );
  sg13g2_a22oi_1 _13326_ (
    .A1(_01382_),
    .A2(_03131_),
    .B1(_03134_),
    .B2(addr_i_9_),
    .Y(_03135_)
  );
  sg13g2_o21ai_1 _13327_ (
    .A1(_00715_),
    .A2(_03130_),
    .B1(_03135_),
    .Y(_03136_)
  );
  sg13g2_nor2_1 _13328_ (
    .A(_00725_),
    .B(_03314_),
    .Y(_03137_)
  );
  sg13g2_o21ai_1 _13329_ (
    .A1(_01436_),
    .A2(_03137_),
    .B1(addr_i_3_),
    .Y(_03138_)
  );
  sg13g2_o21ai_1 _13330_ (
    .A1(_02441_),
    .A2(_03577_),
    .B1(_01244_),
    .Y(_03140_)
  );
  sg13g2_and4_1 _13331_ (
    .A(_01118_),
    .B(_02695_),
    .C(_03138_),
    .D(_03140_),
    .X(_03141_)
  );
  sg13g2_nor2_1 _13332_ (
    .A(addr_i_7_),
    .B(_06010_),
    .Y(_03142_)
  );
  sg13g2_a21oi_1 _13333_ (
    .A1(addr_i_7_),
    .A2(_01168_),
    .B1(addr_i_3_),
    .Y(_03143_)
  );
  sg13g2_nor4_1 _13334_ (
    .A(addr_i_8_),
    .B(_02275_),
    .C(_03142_),
    .D(_03143_),
    .Y(_03144_)
  );
  sg13g2_nor3_1 _13335_ (
    .A(_03136_),
    .B(_03141_),
    .C(_03144_),
    .Y(_03145_)
  );
  sg13g2_a22oi_1 _13336_ (
    .A1(addr_i_9_),
    .A2(_03127_),
    .B1(_03145_),
    .B2(addr_i_10_),
    .Y(_03146_)
  );
  sg13g2_a22oi_1 _13337_ (
    .A1(_03076_),
    .A2(_03100_),
    .B1(addr_i_11_),
    .B2(_03146_),
    .Y(_03147_)
  );
  sg13g2_nand2_1 _13338_ (
    .A(_01125_),
    .B(_00056_),
    .Y(_03148_)
  );
  sg13g2_nor2_1 _13339_ (
    .A(_02196_),
    .B(_08376_),
    .Y(_03149_)
  );
  sg13g2_a22oi_1 _13340_ (
    .A1(addr_i_3_),
    .A2(_03148_),
    .B1(_03149_),
    .B2(_02803_),
    .Y(_03151_)
  );
  sg13g2_and2_1 _13341_ (
    .A(_06496_),
    .B(_01228_),
    .X(_03152_)
  );
  sg13g2_nor3_1 _13342_ (
    .A(addr_i_3_),
    .B(_02053_),
    .C(_03172_),
    .Y(_03153_)
  );
  sg13g2_a21oi_1 _13343_ (
    .A1(addr_i_3_),
    .A2(_03152_),
    .B1(_03153_),
    .Y(_03154_)
  );
  sg13g2_a21oi_1 _13344_ (
    .A1(_03045_),
    .A2(_01747_),
    .B1(_07171_),
    .Y(_03155_)
  );
  sg13g2_o21ai_1 _13345_ (
    .A1(addr_i_2_),
    .A2(_03154_),
    .B1(_03155_),
    .Y(_03156_)
  );
  sg13g2_nor2_1 _13346_ (
    .A(addr_i_4_),
    .B(_03156_),
    .Y(_03157_)
  );
  sg13g2_a21oi_1 _13347_ (
    .A1(addr_i_4_),
    .A2(_00961_),
    .B1(_01507_),
    .Y(_03158_)
  );
  sg13g2_o21ai_1 _13348_ (
    .A1(_00297_),
    .A2(_08144_),
    .B1(_06419_),
    .Y(_03159_)
  );
  sg13g2_o21ai_1 _13349_ (
    .A1(_06154_),
    .A2(_03158_),
    .B1(_03159_),
    .Y(_03160_)
  );
  sg13g2_a21oi_1 _13350_ (
    .A1(addr_i_6_),
    .A2(_03160_),
    .B1(_06695_),
    .Y(_03162_)
  );
  sg13g2_o21ai_1 _13351_ (
    .A1(_03151_),
    .A2(_03157_),
    .B1(_03162_),
    .Y(_03163_)
  );
  sg13g2_a21oi_1 _13352_ (
    .A1(_00441_),
    .A2(_06032_),
    .B1(addr_i_3_),
    .Y(_03164_)
  );
  sg13g2_o21ai_1 _13353_ (
    .A1(_03133_),
    .A2(_03164_),
    .B1(_04052_),
    .Y(_03165_)
  );
  sg13g2_a21oi_1 _13354_ (
    .A1(_00022_),
    .A2(_02746_),
    .B1(_01099_),
    .Y(_03166_)
  );
  sg13g2_buf_1 _13355_ (
    .A(_05899_),
    .X(_03167_)
  );
  sg13g2_a21oi_1 _13356_ (
    .A1(_07724_),
    .A2(_03167_),
    .B1(addr_i_2_),
    .Y(_03168_)
  );
  sg13g2_o21ai_1 _13357_ (
    .A1(_00743_),
    .A2(_03168_),
    .B1(_00799_),
    .Y(_03169_)
  );
  sg13g2_nor2_1 _13358_ (
    .A(addr_i_5_),
    .B(_00447_),
    .Y(_03170_)
  );
  sg13g2_a21oi_1 _13359_ (
    .A1(addr_i_3_),
    .A2(_03061_),
    .B1(_03170_),
    .Y(_03171_)
  );
  sg13g2_a21oi_1 _13360_ (
    .A1(_03169_),
    .A2(_03171_),
    .B1(_00600_),
    .Y(_03173_)
  );
  sg13g2_a21oi_1 _13361_ (
    .A1(_03165_),
    .A2(_03166_),
    .B1(_03173_),
    .Y(_03174_)
  );
  sg13g2_a21oi_1 _13362_ (
    .A1(_03163_),
    .A2(_03174_),
    .B1(_00925_),
    .Y(_03175_)
  );
  sg13g2_nand2_1 _13363_ (
    .A(addr_i_3_),
    .B(_02425_),
    .Y(_03176_)
  );
  sg13g2_nand3_1 _13364_ (
    .A(addr_i_6_),
    .B(_03094_),
    .C(_03176_),
    .Y(_03177_)
  );
  sg13g2_a22oi_1 _13365_ (
    .A1(_00729_),
    .A2(_02742_),
    .B1(_02055_),
    .B2(addr_i_7_),
    .Y(_03178_)
  );
  sg13g2_nand2_1 _13366_ (
    .A(_00210_),
    .B(_00008_),
    .Y(_03179_)
  );
  sg13g2_nand3_1 _13367_ (
    .A(_00262_),
    .B(_02165_),
    .C(_03179_),
    .Y(_03180_)
  );
  sg13g2_nand2_1 _13368_ (
    .A(addr_i_8_),
    .B(_03180_),
    .Y(_03181_)
  );
  sg13g2_nand2_1 _13369_ (
    .A(_08752_),
    .B(_01830_),
    .Y(_03182_)
  );
  sg13g2_a21oi_1 _13370_ (
    .A1(_01287_),
    .A2(_03182_),
    .B1(_00825_),
    .Y(_03184_)
  );
  sg13g2_a22oi_1 _13371_ (
    .A1(_03177_),
    .A2(_03178_),
    .B1(_03181_),
    .B2(_03184_),
    .Y(_03185_)
  );
  sg13g2_nor2_1 _13372_ (
    .A(_04075_),
    .B(_01724_),
    .Y(_03186_)
  );
  sg13g2_a22oi_1 _13373_ (
    .A1(addr_i_3_),
    .A2(_02410_),
    .B1(_03186_),
    .B2(_02213_),
    .Y(_03187_)
  );
  sg13g2_nor2_1 _13374_ (
    .A(_03765_),
    .B(_05943_),
    .Y(_03188_)
  );
  sg13g2_nand2_1 _13375_ (
    .A(addr_i_4_),
    .B(_03188_),
    .Y(_03189_)
  );
  sg13g2_nor2_1 _13376_ (
    .A(addr_i_5_),
    .B(_00208_),
    .Y(_03190_)
  );
  sg13g2_nand2_1 _13377_ (
    .A(_01113_),
    .B(_03190_),
    .Y(_03191_)
  );
  sg13g2_a21oi_1 _13378_ (
    .A1(_03189_),
    .A2(_03191_),
    .B1(_00021_),
    .Y(_03192_)
  );
  sg13g2_or3_1 _13379_ (
    .A(addr_i_8_),
    .B(_03187_),
    .C(_03192_),
    .X(_03193_)
  );
  sg13g2_nor2_1 _13380_ (
    .A(_06176_),
    .B(_08288_),
    .Y(_03195_)
  );
  sg13g2_nor3_1 _13381_ (
    .A(addr_i_3_),
    .B(_00597_),
    .C(_00426_),
    .Y(_03196_)
  );
  sg13g2_a22oi_1 _13382_ (
    .A1(addr_i_3_),
    .A2(_03195_),
    .B1(_03196_),
    .B2(addr_i_4_),
    .Y(_03197_)
  );
  sg13g2_a22oi_1 _13383_ (
    .A1(_01019_),
    .A2(_02008_),
    .B1(_03197_),
    .B2(_05822_),
    .Y(_03198_)
  );
  sg13g2_o21ai_1 _13384_ (
    .A1(_03193_),
    .A2(_03198_),
    .B1(_01174_),
    .Y(_03199_)
  );
  sg13g2_o21ai_1 _13385_ (
    .A1(_04151_),
    .A2(_03110_),
    .B1(_00034_),
    .Y(_03200_)
  );
  sg13g2_nand2_1 _13386_ (
    .A(addr_i_2_),
    .B(_03200_),
    .Y(_03201_)
  );
  sg13g2_o21ai_1 _13387_ (
    .A1(_06497_),
    .A2(_00885_),
    .B1(addr_i_4_),
    .Y(_03202_)
  );
  sg13g2_nand2_1 _13388_ (
    .A(_05070_),
    .B(_02952_),
    .Y(_03203_)
  );
  sg13g2_a22oi_1 _13389_ (
    .A1(_00375_),
    .A2(_09510_),
    .B1(_03203_),
    .B2(addr_i_10_),
    .Y(_03204_)
  );
  sg13g2_nand3_1 _13390_ (
    .A(_03201_),
    .B(_03202_),
    .C(_03204_),
    .Y(_03206_)
  );
  sg13g2_and2_1 _13391_ (
    .A(addr_i_11_),
    .B(_03206_),
    .X(_03207_)
  );
  sg13g2_o21ai_1 _13392_ (
    .A1(_03185_),
    .A2(_03199_),
    .B1(_03207_),
    .Y(_03208_)
  );
  sg13g2_nor2_1 _13393_ (
    .A(addr_i_5_),
    .B(_01254_),
    .Y(_03209_)
  );
  sg13g2_nand2_1 _13394_ (
    .A(_05546_),
    .B(_00671_),
    .Y(_03210_)
  );
  sg13g2_a22oi_1 _13395_ (
    .A1(_02105_),
    .A2(_03210_),
    .B1(_00376_),
    .B2(_02063_),
    .Y(_03211_)
  );
  sg13g2_nand2_1 _13396_ (
    .A(addr_i_3_),
    .B(_01765_),
    .Y(_03212_)
  );
  sg13g2_o21ai_1 _13397_ (
    .A1(_03209_),
    .A2(_03211_),
    .B1(_03212_),
    .Y(_03213_)
  );
  sg13g2_a21oi_1 _13398_ (
    .A1(addr_i_7_),
    .A2(_03213_),
    .B1(_00367_),
    .Y(_03214_)
  );
  sg13g2_o21ai_1 _13399_ (
    .A1(_00292_),
    .A2(_00990_),
    .B1(addr_i_4_),
    .Y(_03215_)
  );
  sg13g2_a21oi_1 _13400_ (
    .A1(addr_i_2_),
    .A2(_08796_),
    .B1(addr_i_4_),
    .Y(_03217_)
  );
  sg13g2_o21ai_1 _13401_ (
    .A1(_09494_),
    .A2(_03217_),
    .B1(addr_i_7_),
    .Y(_03218_)
  );
  sg13g2_nand4_1 _13402_ (
    .A(addr_i_3_),
    .B(_00405_),
    .C(_03215_),
    .D(_03218_),
    .Y(_03219_)
  );
  sg13g2_o21ai_1 _13403_ (
    .A1(_02238_),
    .A2(_06563_),
    .B1(addr_i_4_),
    .Y(_03220_)
  );
  sg13g2_nor3_1 _13404_ (
    .A(addr_i_4_),
    .B(addr_i_6_),
    .C(_00165_),
    .Y(_03221_)
  );
  sg13g2_o21ai_1 _13405_ (
    .A1(_01972_),
    .A2(_03221_),
    .B1(addr_i_2_),
    .Y(_03222_)
  );
  sg13g2_nand4_1 _13406_ (
    .A(_00701_),
    .B(_00677_),
    .C(_03220_),
    .D(_03222_),
    .Y(_03223_)
  );
  sg13g2_a221oi_1 _13407_ (
    .A1(_00292_),
    .A2(_00574_),
    .B1(_03219_),
    .B2(_03223_),
    .C1(addr_i_8_),
    .Y(_03224_)
  );
  sg13g2_nor3_1 _13408_ (
    .A(_00774_),
    .B(_03214_),
    .C(_03224_),
    .Y(_03225_)
  );
  sg13g2_buf_1 _13409_ (
    .A(_00785_),
    .X(_03226_)
  );
  sg13g2_nand2_1 _13410_ (
    .A(_00339_),
    .B(_03226_),
    .Y(_03228_)
  );
  sg13g2_nand2_1 _13411_ (
    .A(_00770_),
    .B(_08464_),
    .Y(_03229_)
  );
  sg13g2_nor2_1 _13412_ (
    .A(_00644_),
    .B(_03229_),
    .Y(_03230_)
  );
  sg13g2_a21oi_1 _13413_ (
    .A1(_00467_),
    .A2(_00148_),
    .B1(addr_i_2_),
    .Y(_03231_)
  );
  sg13g2_a22oi_1 _13414_ (
    .A1(addr_i_3_),
    .A2(_03228_),
    .B1(_03230_),
    .B2(_03231_),
    .Y(_03232_)
  );
  sg13g2_nor2_1 _13415_ (
    .A(addr_i_6_),
    .B(_05346_),
    .Y(_03233_)
  );
  sg13g2_o21ai_1 _13416_ (
    .A1(addr_i_3_),
    .A2(_03233_),
    .B1(_00477_),
    .Y(_03234_)
  );
  sg13g2_nand2_1 _13417_ (
    .A(_05036_),
    .B(_05379_),
    .Y(_03235_)
  );
  sg13g2_a21oi_1 _13418_ (
    .A1(_09478_),
    .A2(_03235_),
    .B1(addr_i_4_),
    .Y(_03236_)
  );
  sg13g2_a22oi_1 _13419_ (
    .A1(addr_i_4_),
    .A2(_03234_),
    .B1(_03236_),
    .B2(_00474_),
    .Y(_03237_)
  );
  sg13g2_nand2_1 _13420_ (
    .A(addr_i_7_),
    .B(_03237_),
    .Y(_03239_)
  );
  sg13g2_o21ai_1 _13421_ (
    .A1(addr_i_7_),
    .A2(_03232_),
    .B1(_03239_),
    .Y(_03240_)
  );
  sg13g2_xnor2_1 _13422_ (
    .A(addr_i_3_),
    .B(_05501_),
    .Y(_03241_)
  );
  sg13g2_o21ai_1 _13423_ (
    .A1(_00051_),
    .A2(_03241_),
    .B1(addr_i_8_),
    .Y(_03242_)
  );
  sg13g2_nor2_1 _13424_ (
    .A(_04041_),
    .B(_09497_),
    .Y(_03243_)
  );
  sg13g2_o21ai_1 _13425_ (
    .A1(addr_i_3_),
    .A2(_03243_),
    .B1(_00704_),
    .Y(_03244_)
  );
  sg13g2_buf_1 _13426_ (
    .A(_00890_),
    .X(_03245_)
  );
  sg13g2_o21ai_1 _13427_ (
    .A1(_03245_),
    .A2(_00632_),
    .B1(addr_i_4_),
    .Y(_03246_)
  );
  sg13g2_a21oi_1 _13428_ (
    .A1(_09260_),
    .A2(_03246_),
    .B1(_01169_),
    .Y(_03247_)
  );
  sg13g2_nand2_1 _13429_ (
    .A(addr_i_3_),
    .B(_07027_),
    .Y(_03248_)
  );
  sg13g2_nand2_1 _13430_ (
    .A(_00413_),
    .B(_08221_),
    .Y(_03250_)
  );
  sg13g2_nand2_1 _13431_ (
    .A(_07503_),
    .B(_03250_),
    .Y(_03251_)
  );
  sg13g2_a21oi_1 _13432_ (
    .A1(_03248_),
    .A2(_03251_),
    .B1(addr_i_5_),
    .Y(_03252_)
  );
  sg13g2_a22oi_1 _13433_ (
    .A1(_01475_),
    .A2(_03244_),
    .B1(_03247_),
    .B2(_03252_),
    .Y(_03253_)
  );
  sg13g2_nor2_1 _13434_ (
    .A(_03242_),
    .B(_03253_),
    .Y(_03254_)
  );
  sg13g2_a22oi_1 _13435_ (
    .A1(_00114_),
    .A2(_03240_),
    .B1(_03254_),
    .B2(_01452_),
    .Y(_03255_)
  );
  sg13g2_nor4_1 _13436_ (
    .A(_03175_),
    .B(_03208_),
    .C(_03225_),
    .D(_03255_),
    .Y(_03256_)
  );
  sg13g2_or3_1 _13437_ (
    .A(addr_i_12_),
    .B(_03147_),
    .C(_03256_),
    .X(_03257_)
  );
  sg13g2_o21ai_1 _13438_ (
    .A1(_03028_),
    .A2(_03057_),
    .B1(_03257_),
    .Y(data_o_17_)
  );
  sg13g2_nand2_1 _13439_ (
    .A(_08044_),
    .B(_03110_),
    .Y(_03258_)
  );
  sg13g2_buf_1 _13440_ (
    .A(_01674_),
    .X(_03260_)
  );
  sg13g2_nor2_1 _13441_ (
    .A(_03260_),
    .B(_02772_),
    .Y(_03261_)
  );
  sg13g2_nor2_1 _13442_ (
    .A(addr_i_5_),
    .B(_07636_),
    .Y(_03262_)
  );
  sg13g2_buf_1 _13443_ (
    .A(_03776_),
    .X(_03263_)
  );
  sg13g2_a21oi_1 _13444_ (
    .A1(_02528_),
    .A2(_02683_),
    .B1(_03263_),
    .Y(_03264_)
  );
  sg13g2_a22oi_1 _13445_ (
    .A1(_08399_),
    .A2(_03262_),
    .B1(_03264_),
    .B2(addr_i_3_),
    .Y(_03265_)
  );
  sg13g2_a22oi_1 _13446_ (
    .A1(_03258_),
    .A2(_03261_),
    .B1(_03265_),
    .B2(_03062_),
    .Y(_03266_)
  );
  sg13g2_nor2_1 _13447_ (
    .A(addr_i_3_),
    .B(_04726_),
    .Y(_03267_)
  );
  sg13g2_a21oi_1 _13448_ (
    .A1(addr_i_3_),
    .A2(_01057_),
    .B1(_03267_),
    .Y(_03268_)
  );
  sg13g2_or2_1 _13449_ (
    .A(_05999_),
    .B(_01654_),
    .X(_03269_)
  );
  sg13g2_a22oi_1 _13450_ (
    .A1(addr_i_2_),
    .A2(_03269_),
    .B1(_01031_),
    .B2(_00860_),
    .Y(_03271_)
  );
  sg13g2_o21ai_1 _13451_ (
    .A1(addr_i_5_),
    .A2(_03268_),
    .B1(_03271_),
    .Y(_03272_)
  );
  sg13g2_nand2_1 _13452_ (
    .A(_00072_),
    .B(_04162_),
    .Y(_03273_)
  );
  sg13g2_a21oi_1 _13453_ (
    .A1(_00747_),
    .A2(_03273_),
    .B1(_00492_),
    .Y(_03274_)
  );
  sg13g2_o21ai_1 _13454_ (
    .A1(_08310_),
    .A2(_03274_),
    .B1(addr_i_8_),
    .Y(_03275_)
  );
  sg13g2_a22oi_1 _13455_ (
    .A1(_00697_),
    .A2(_01125_),
    .B1(_00125_),
    .B2(_07514_),
    .Y(_03276_)
  );
  sg13g2_a22oi_1 _13456_ (
    .A1(_09205_),
    .A2(_01354_),
    .B1(addr_i_4_),
    .B2(_07514_),
    .Y(_03277_)
  );
  sg13g2_a221oi_1 _13457_ (
    .A1(addr_i_3_),
    .A2(_01001_),
    .B1(_02380_),
    .B2(_00381_),
    .C1(_07945_),
    .Y(_03278_)
  );
  sg13g2_nor4_1 _13458_ (
    .A(_00385_),
    .B(_03276_),
    .C(_03277_),
    .D(_03278_),
    .Y(_03279_)
  );
  sg13g2_nand3_1 _13459_ (
    .A(_03272_),
    .B(_03275_),
    .C(_03279_),
    .Y(_03280_)
  );
  sg13g2_a21oi_1 _13460_ (
    .A1(_00549_),
    .A2(_01745_),
    .B1(_01888_),
    .Y(_03282_)
  );
  sg13g2_nor2_1 _13461_ (
    .A(_01592_),
    .B(_01652_),
    .Y(_03283_)
  );
  sg13g2_nor2_1 _13462_ (
    .A(_02371_),
    .B(_02196_),
    .Y(_03284_)
  );
  sg13g2_o21ai_1 _13463_ (
    .A1(_03283_),
    .A2(_03284_),
    .B1(addr_i_4_),
    .Y(_03285_)
  );
  sg13g2_o21ai_1 _13464_ (
    .A1(addr_i_5_),
    .A2(_03282_),
    .B1(_03285_),
    .Y(_03286_)
  );
  sg13g2_nor2_1 _13465_ (
    .A(_03820_),
    .B(_00034_),
    .Y(_03287_)
  );
  sg13g2_buf_1 _13466_ (
    .A(_05379_),
    .X(_03288_)
  );
  sg13g2_nand2_1 _13467_ (
    .A(_00078_),
    .B(_02254_),
    .Y(_03289_)
  );
  sg13g2_a21oi_1 _13468_ (
    .A1(_06851_),
    .A2(_00975_),
    .B1(addr_i_3_),
    .Y(_03290_)
  );
  sg13g2_a21oi_1 _13469_ (
    .A1(_03288_),
    .A2(_03289_),
    .B1(_03290_),
    .Y(_03291_)
  );
  sg13g2_a21oi_1 _13470_ (
    .A1(_02546_),
    .A2(_03291_),
    .B1(addr_i_5_),
    .Y(_03293_)
  );
  sg13g2_a221oi_1 _13471_ (
    .A1(addr_i_6_),
    .A2(_03286_),
    .B1(_03287_),
    .B2(_03045_),
    .C1(_03293_),
    .Y(_03294_)
  );
  sg13g2_a21oi_1 _13472_ (
    .A1(_09205_),
    .A2(_01060_),
    .B1(_01308_),
    .Y(_03295_)
  );
  sg13g2_o21ai_1 _13473_ (
    .A1(_02772_),
    .A2(_03295_),
    .B1(addr_i_4_),
    .Y(_03296_)
  );
  sg13g2_o21ai_1 _13474_ (
    .A1(addr_i_3_),
    .A2(_03112_),
    .B1(_00582_),
    .Y(_03297_)
  );
  sg13g2_a22oi_1 _13475_ (
    .A1(_02277_),
    .A2(_03297_),
    .B1(_00945_),
    .B2(_03227_),
    .Y(_03298_)
  );
  sg13g2_nand2_1 _13476_ (
    .A(_09393_),
    .B(_09404_),
    .Y(_03299_)
  );
  sg13g2_nor2_1 _13477_ (
    .A(addr_i_3_),
    .B(_03299_),
    .Y(_03300_)
  );
  sg13g2_a22oi_1 _13478_ (
    .A1(addr_i_3_),
    .A2(_04727_),
    .B1(_03300_),
    .B2(_01131_),
    .Y(_03301_)
  );
  sg13g2_a22oi_1 _13479_ (
    .A1(_00990_),
    .A2(_00861_),
    .B1(_09459_),
    .B2(addr_i_4_),
    .Y(_03302_)
  );
  sg13g2_nor3_1 _13480_ (
    .A(_01285_),
    .B(_03301_),
    .C(_03302_),
    .Y(_03304_)
  );
  sg13g2_a22oi_1 _13481_ (
    .A1(_03296_),
    .A2(_03298_),
    .B1(addr_i_9_),
    .B2(_03304_),
    .Y(_03305_)
  );
  sg13g2_o21ai_1 _13482_ (
    .A1(addr_i_8_),
    .A2(_03294_),
    .B1(_03305_),
    .Y(_03306_)
  );
  sg13g2_o21ai_1 _13483_ (
    .A1(_03266_),
    .A2(_03280_),
    .B1(_03306_),
    .Y(_03307_)
  );
  sg13g2_nor2_1 _13484_ (
    .A(_01384_),
    .B(_08941_),
    .Y(_03308_)
  );
  sg13g2_o21ai_1 _13485_ (
    .A1(_03308_),
    .A2(_01540_),
    .B1(addr_i_6_),
    .Y(_03309_)
  );
  sg13g2_a21oi_1 _13486_ (
    .A1(_06862_),
    .A2(_03864_),
    .B1(_03776_),
    .Y(_03310_)
  );
  sg13g2_a21oi_1 _13487_ (
    .A1(_03288_),
    .A2(_02536_),
    .B1(_03310_),
    .Y(_03311_)
  );
  sg13g2_nand4_1 _13488_ (
    .A(_00351_),
    .B(_07569_),
    .C(_03309_),
    .D(_03311_),
    .Y(_03312_)
  );
  sg13g2_a21oi_1 _13489_ (
    .A1(_06884_),
    .A2(_01406_),
    .B1(addr_i_3_),
    .Y(_03313_)
  );
  sg13g2_o21ai_1 _13490_ (
    .A1(_01986_),
    .A2(_03313_),
    .B1(addr_i_4_),
    .Y(_03315_)
  );
  sg13g2_o21ai_1 _13491_ (
    .A1(_00282_),
    .A2(_01478_),
    .B1(_08155_),
    .Y(_03316_)
  );
  sg13g2_nand4_1 _13492_ (
    .A(addr_i_7_),
    .B(_00470_),
    .C(_03315_),
    .D(_03316_),
    .Y(_03317_)
  );
  sg13g2_nand2_1 _13493_ (
    .A(_03312_),
    .B(_03317_),
    .Y(_03318_)
  );
  sg13g2_a21oi_1 _13494_ (
    .A1(addr_i_3_),
    .A2(_01572_),
    .B1(_02639_),
    .Y(_03319_)
  );
  sg13g2_o21ai_1 _13495_ (
    .A1(_03032_),
    .A2(_01281_),
    .B1(addr_i_7_),
    .Y(_03320_)
  );
  sg13g2_a21o_1 _13496_ (
    .A1(_00050_),
    .A2(_03320_),
    .B1(addr_i_2_),
    .X(_03321_)
  );
  sg13g2_o21ai_1 _13497_ (
    .A1(_00949_),
    .A2(_03319_),
    .B1(_03321_),
    .Y(_03322_)
  );
  sg13g2_nor2_1 _13498_ (
    .A(_09493_),
    .B(_00252_),
    .Y(_03323_)
  );
  sg13g2_nand2_1 _13499_ (
    .A(_05324_),
    .B(_07237_),
    .Y(_03324_)
  );
  sg13g2_a21oi_1 _13500_ (
    .A1(_03323_),
    .A2(_03324_),
    .B1(_08332_),
    .Y(_03326_)
  );
  sg13g2_a21oi_1 _13501_ (
    .A1(addr_i_5_),
    .A2(_00408_),
    .B1(_03358_),
    .Y(_03327_)
  );
  sg13g2_a22oi_1 _13502_ (
    .A1(_01881_),
    .A2(_02976_),
    .B1(_03326_),
    .B2(_03327_),
    .Y(_03328_)
  );
  sg13g2_nor2_1 _13503_ (
    .A(_04052_),
    .B(_03328_),
    .Y(_03329_)
  );
  sg13g2_o21ai_1 _13504_ (
    .A1(_03322_),
    .A2(_03329_),
    .B1(addr_i_8_),
    .Y(_03330_)
  );
  sg13g2_o21ai_1 _13505_ (
    .A1(addr_i_8_),
    .A2(_03318_),
    .B1(_03330_),
    .Y(_03331_)
  );
  sg13g2_o21ai_1 _13506_ (
    .A1(_09494_),
    .A2(_09502_),
    .B1(addr_i_3_),
    .Y(_03332_)
  );
  sg13g2_nand2_1 _13507_ (
    .A(_01967_),
    .B(_03332_),
    .Y(_03333_)
  );
  sg13g2_o21ai_1 _13508_ (
    .A1(_02064_),
    .A2(_01450_),
    .B1(_03853_),
    .Y(_03334_)
  );
  sg13g2_nand3_1 _13509_ (
    .A(addr_i_2_),
    .B(_00077_),
    .C(_03334_),
    .Y(_03335_)
  );
  sg13g2_o21ai_1 _13510_ (
    .A1(addr_i_2_),
    .A2(_03333_),
    .B1(_03335_),
    .Y(_03337_)
  );
  sg13g2_o21ai_1 _13511_ (
    .A1(_00414_),
    .A2(_00258_),
    .B1(_01073_),
    .Y(_03338_)
  );
  sg13g2_nand2_1 _13512_ (
    .A(_07282_),
    .B(_00405_),
    .Y(_03339_)
  );
  sg13g2_nand2_1 _13513_ (
    .A(_01585_),
    .B(_05501_),
    .Y(_03340_)
  );
  sg13g2_a21oi_1 _13514_ (
    .A1(_02898_),
    .A2(_03340_),
    .B1(addr_i_3_),
    .Y(_03341_)
  );
  sg13g2_a22oi_1 _13515_ (
    .A1(addr_i_5_),
    .A2(_03338_),
    .B1(_03339_),
    .B2(_03341_),
    .Y(_03342_)
  );
  sg13g2_a221oi_1 _13516_ (
    .A1(addr_i_4_),
    .A2(_01319_),
    .B1(_00110_),
    .B2(_00915_),
    .C1(_00534_),
    .Y(_03343_)
  );
  sg13g2_a221oi_1 _13517_ (
    .A1(addr_i_3_),
    .A2(_05280_),
    .B1(_07458_),
    .B2(_02426_),
    .C1(_05999_),
    .Y(_03344_)
  );
  sg13g2_o21ai_1 _13518_ (
    .A1(addr_i_3_),
    .A2(_03343_),
    .B1(_03344_),
    .Y(_03345_)
  );
  sg13g2_nand2_1 _13519_ (
    .A(_01159_),
    .B(_00238_),
    .Y(_03346_)
  );
  sg13g2_buf_1 _13520_ (
    .A(_01943_),
    .X(_03348_)
  );
  sg13g2_o21ai_1 _13521_ (
    .A1(addr_i_6_),
    .A2(_00292_),
    .B1(_03348_),
    .Y(_03349_)
  );
  sg13g2_nand2_1 _13522_ (
    .A(_05236_),
    .B(_01652_),
    .Y(_03350_)
  );
  sg13g2_nand3_1 _13523_ (
    .A(_03346_),
    .B(_03349_),
    .C(_03350_),
    .Y(_03351_)
  );
  sg13g2_o21ai_1 _13524_ (
    .A1(addr_i_2_),
    .A2(_02150_),
    .B1(addr_i_8_),
    .Y(_03352_)
  );
  sg13g2_a221oi_1 _13525_ (
    .A1(addr_i_2_),
    .A2(_03345_),
    .B1(_03351_),
    .B2(_08399_),
    .C1(_03352_),
    .Y(_03353_)
  );
  sg13g2_a22oi_1 _13526_ (
    .A1(_03337_),
    .A2(_03342_),
    .B1(_03353_),
    .B2(addr_i_9_),
    .Y(_03354_)
  );
  sg13g2_a22oi_1 _13527_ (
    .A1(addr_i_9_),
    .A2(_03331_),
    .B1(_03354_),
    .B2(addr_i_10_),
    .Y(_03355_)
  );
  sg13g2_a21oi_1 _13528_ (
    .A1(addr_i_10_),
    .A2(_03307_),
    .B1(_03355_),
    .Y(_03356_)
  );
  sg13g2_nand4_1 _13529_ (
    .A(_09487_),
    .B(_05490_),
    .C(_02604_),
    .D(_01097_),
    .Y(_03357_)
  );
  sg13g2_inv_1 _13530_ (
    .A(_01398_),
    .Y(_03359_)
  );
  sg13g2_a21oi_1 _13531_ (
    .A1(_09105_),
    .A2(_06873_),
    .B1(addr_i_3_),
    .Y(_03360_)
  );
  sg13g2_nor2_1 _13532_ (
    .A(_00317_),
    .B(_01611_),
    .Y(_03361_)
  );
  sg13g2_o21ai_1 _13533_ (
    .A1(_03359_),
    .A2(_03360_),
    .B1(_03361_),
    .Y(_03362_)
  );
  sg13g2_nand3_1 _13534_ (
    .A(addr_i_10_),
    .B(_03357_),
    .C(_03362_),
    .Y(_03363_)
  );
  sg13g2_nand2_1 _13535_ (
    .A(_00520_),
    .B(_07790_),
    .Y(_03364_)
  );
  sg13g2_o21ai_1 _13536_ (
    .A1(_00838_),
    .A2(_01007_),
    .B1(_01368_),
    .Y(_03365_)
  );
  sg13g2_a221oi_1 _13537_ (
    .A1(_00500_),
    .A2(_03364_),
    .B1(_03365_),
    .B2(_08011_),
    .C1(addr_i_7_),
    .Y(_03366_)
  );
  sg13g2_a21oi_1 _13538_ (
    .A1(_02513_),
    .A2(_02529_),
    .B1(_08266_),
    .Y(_03367_)
  );
  sg13g2_o21ai_1 _13539_ (
    .A1(_09105_),
    .A2(_05114_),
    .B1(addr_i_7_),
    .Y(_03368_)
  );
  sg13g2_o21ai_1 _13540_ (
    .A1(_03367_),
    .A2(_03368_),
    .B1(_00423_),
    .Y(_03370_)
  );
  sg13g2_nand2_1 _13541_ (
    .A(_06220_),
    .B(_07900_),
    .Y(_03371_)
  );
  sg13g2_nand2_1 _13542_ (
    .A(_00749_),
    .B(_03371_),
    .Y(_03372_)
  );
  sg13g2_a21oi_1 _13543_ (
    .A1(_00820_),
    .A2(_00603_),
    .B1(addr_i_4_),
    .Y(_03373_)
  );
  sg13g2_nor2_1 _13544_ (
    .A(_05811_),
    .B(_01610_),
    .Y(_03374_)
  );
  sg13g2_o21ai_1 _13545_ (
    .A1(_03372_),
    .A2(_03373_),
    .B1(_03374_),
    .Y(_03375_)
  );
  sg13g2_o21ai_1 _13546_ (
    .A1(_03366_),
    .A2(_03370_),
    .B1(_03375_),
    .Y(_03376_)
  );
  sg13g2_a21oi_1 _13547_ (
    .A1(_01262_),
    .A2(_00594_),
    .B1(_01732_),
    .Y(_03377_)
  );
  sg13g2_o21ai_1 _13548_ (
    .A1(_04284_),
    .A2(_06939_),
    .B1(addr_i_2_),
    .Y(_03378_)
  );
  sg13g2_o21ai_1 _13549_ (
    .A1(_07193_),
    .A2(_00209_),
    .B1(_00956_),
    .Y(_03379_)
  );
  sg13g2_nand3_1 _13550_ (
    .A(_01734_),
    .B(_03378_),
    .C(_03379_),
    .Y(_03381_)
  );
  sg13g2_a21oi_1 _13551_ (
    .A1(addr_i_7_),
    .A2(_06077_),
    .B1(_04362_),
    .Y(_03382_)
  );
  sg13g2_nor2_1 _13552_ (
    .A(_02134_),
    .B(_03382_),
    .Y(_03383_)
  );
  sg13g2_nor2_1 _13553_ (
    .A(_05003_),
    .B(_09506_),
    .Y(_03384_)
  );
  sg13g2_o21ai_1 _13554_ (
    .A1(_03383_),
    .A2(_03384_),
    .B1(addr_i_3_),
    .Y(_03385_)
  );
  sg13g2_o21ai_1 _13555_ (
    .A1(addr_i_3_),
    .A2(_03381_),
    .B1(_03385_),
    .Y(_03386_)
  );
  sg13g2_o21ai_1 _13556_ (
    .A1(addr_i_4_),
    .A2(_03377_),
    .B1(_03386_),
    .Y(_03387_)
  );
  sg13g2_nand2_1 _13557_ (
    .A(_00554_),
    .B(_01212_),
    .Y(_03388_)
  );
  sg13g2_a21oi_1 _13558_ (
    .A1(_00103_),
    .A2(_03388_),
    .B1(_08431_),
    .Y(_03389_)
  );
  sg13g2_nand2b_1 _13559_ (
    .A_N(_01016_),
    .B(_01857_),
    .Y(_03390_)
  );
  sg13g2_nor3_1 _13560_ (
    .A(addr_i_8_),
    .B(_03389_),
    .C(_03390_),
    .Y(_03392_)
  );
  sg13g2_nand2_1 _13561_ (
    .A(_01672_),
    .B(_02012_),
    .Y(_03393_)
  );
  sg13g2_a21oi_1 _13562_ (
    .A1(_00477_),
    .A2(_03248_),
    .B1(_00554_),
    .Y(_03394_)
  );
  sg13g2_a22oi_1 _13563_ (
    .A1(_00190_),
    .A2(_03393_),
    .B1(_03394_),
    .B2(_00247_),
    .Y(_03395_)
  );
  sg13g2_nand2b_1 _13564_ (
    .A_N(_03395_),
    .B(addr_i_5_),
    .Y(_03396_)
  );
  sg13g2_a221oi_1 _13565_ (
    .A1(addr_i_8_),
    .A2(_03387_),
    .B1(_03392_),
    .B2(_03396_),
    .C1(_00396_),
    .Y(_03397_)
  );
  sg13g2_nor3_1 _13566_ (
    .A(_03363_),
    .B(_03376_),
    .C(_03397_),
    .Y(_03398_)
  );
  sg13g2_nor2_1 _13567_ (
    .A(_00065_),
    .B(_02312_),
    .Y(_03399_)
  );
  sg13g2_a21oi_1 _13568_ (
    .A1(addr_i_7_),
    .A2(_03545_),
    .B1(_03399_),
    .Y(_03400_)
  );
  sg13g2_nor2_1 _13569_ (
    .A(_03446_),
    .B(_05390_),
    .Y(_03401_)
  );
  sg13g2_a21oi_1 _13570_ (
    .A1(_09486_),
    .A2(_03401_),
    .B1(_00029_),
    .Y(_03403_)
  );
  sg13g2_o21ai_1 _13571_ (
    .A1(addr_i_4_),
    .A2(_03400_),
    .B1(_03403_),
    .Y(_03404_)
  );
  sg13g2_o21ai_1 _13572_ (
    .A1(addr_i_7_),
    .A2(_05424_),
    .B1(addr_i_2_),
    .Y(_03405_)
  );
  sg13g2_nand2_1 _13573_ (
    .A(_06784_),
    .B(_03405_),
    .Y(_03406_)
  );
  sg13g2_a22oi_1 _13574_ (
    .A1(_00052_),
    .A2(_00516_),
    .B1(addr_i_4_),
    .B2(addr_i_2_),
    .Y(_03407_)
  );
  sg13g2_a22oi_1 _13575_ (
    .A1(addr_i_4_),
    .A2(_03406_),
    .B1(_03407_),
    .B2(_00898_),
    .Y(_03408_)
  );
  sg13g2_nor2_1 _13576_ (
    .A(addr_i_3_),
    .B(_03408_),
    .Y(_03409_)
  );
  sg13g2_nand2_1 _13577_ (
    .A(addr_i_8_),
    .B(_01586_),
    .Y(_03410_)
  );
  sg13g2_a22oi_1 _13578_ (
    .A1(addr_i_3_),
    .A2(_03404_),
    .B1(_03409_),
    .B2(_03410_),
    .Y(_03411_)
  );
  sg13g2_or2_1 _13579_ (
    .A(_00257_),
    .B(_02123_),
    .X(_03412_)
  );
  sg13g2_nor3_1 _13580_ (
    .A(_02976_),
    .B(_00034_),
    .C(_03245_),
    .Y(_03414_)
  );
  sg13g2_a22oi_1 _13581_ (
    .A1(addr_i_4_),
    .A2(_03412_),
    .B1(_03414_),
    .B2(addr_i_5_),
    .Y(_03415_)
  );
  sg13g2_nor2_1 _13582_ (
    .A(_00435_),
    .B(_08453_),
    .Y(_03416_)
  );
  sg13g2_a22oi_1 _13583_ (
    .A1(_00157_),
    .A2(_00098_),
    .B1(_03416_),
    .B2(_03263_),
    .Y(_03417_)
  );
  sg13g2_o21ai_1 _13584_ (
    .A1(_03415_),
    .A2(_03417_),
    .B1(_01043_),
    .Y(_03418_)
  );
  sg13g2_nor2b_1 _13585_ (
    .A(_03411_),
    .B_N(_03418_),
    .Y(_03419_)
  );
  sg13g2_nand2_1 _13586_ (
    .A(_08044_),
    .B(_01680_),
    .Y(_03420_)
  );
  sg13g2_nand2_1 _13587_ (
    .A(_02213_),
    .B(_03420_),
    .Y(_03421_)
  );
  sg13g2_a22oi_1 _13588_ (
    .A1(_00190_),
    .A2(_03421_),
    .B1(_00096_),
    .B2(addr_i_5_),
    .Y(_03422_)
  );
  sg13g2_nand2_1 _13589_ (
    .A(_01948_),
    .B(_07116_),
    .Y(_03423_)
  );
  sg13g2_a221oi_1 _13590_ (
    .A1(_01159_),
    .A2(_01445_),
    .B1(_03423_),
    .B2(addr_i_3_),
    .C1(_08708_),
    .Y(_03425_)
  );
  sg13g2_or2_1 _13591_ (
    .A(_03422_),
    .B(_03425_),
    .X(_03426_)
  );
  sg13g2_or2_1 _13592_ (
    .A(_08575_),
    .B(_02180_),
    .X(_03427_)
  );
  sg13g2_nand2_1 _13593_ (
    .A(_00483_),
    .B(_00173_),
    .Y(_03428_)
  );
  sg13g2_nand3_1 _13594_ (
    .A(_00704_),
    .B(_01462_),
    .C(_03428_),
    .Y(_03429_)
  );
  sg13g2_a221oi_1 _13595_ (
    .A1(_00402_),
    .A2(_03427_),
    .B1(_03429_),
    .B2(_01320_),
    .C1(addr_i_8_),
    .Y(_03430_)
  );
  sg13g2_buf_1 _13596_ (
    .A(_00914_),
    .X(_03431_)
  );
  sg13g2_o21ai_1 _13597_ (
    .A1(addr_i_4_),
    .A2(_01508_),
    .B1(_03431_),
    .Y(_03432_)
  );
  sg13g2_nor2_1 _13598_ (
    .A(_02283_),
    .B(_00718_),
    .Y(_03433_)
  );
  sg13g2_a21oi_1 _13599_ (
    .A1(_01262_),
    .A2(_02012_),
    .B1(_03433_),
    .Y(_03434_)
  );
  sg13g2_o21ai_1 _13600_ (
    .A1(_08653_),
    .A2(_00087_),
    .B1(addr_i_4_),
    .Y(_03436_)
  );
  sg13g2_nand3_1 _13601_ (
    .A(addr_i_8_),
    .B(_03434_),
    .C(_03436_),
    .Y(_03437_)
  );
  sg13g2_o21ai_1 _13602_ (
    .A1(_06927_),
    .A2(_02322_),
    .B1(addr_i_3_),
    .Y(_03438_)
  );
  sg13g2_o21ai_1 _13603_ (
    .A1(_06806_),
    .A2(_03720_),
    .B1(_01191_),
    .Y(_03439_)
  );
  sg13g2_a21oi_1 _13604_ (
    .A1(_03438_),
    .A2(_03439_),
    .B1(_00146_),
    .Y(_03440_)
  );
  sg13g2_a22oi_1 _13605_ (
    .A1(_01519_),
    .A2(_03432_),
    .B1(_03437_),
    .B2(_03440_),
    .Y(_03441_)
  );
  sg13g2_a22oi_1 _13606_ (
    .A1(_03426_),
    .A2(_03430_),
    .B1(_03441_),
    .B2(_00243_),
    .Y(_03442_)
  );
  sg13g2_a22oi_1 _13607_ (
    .A1(_00397_),
    .A2(_03419_),
    .B1(_03442_),
    .B2(addr_i_10_),
    .Y(_03443_)
  );
  sg13g2_nor2_1 _13608_ (
    .A(_03398_),
    .B(_03443_),
    .Y(_03444_)
  );
  sg13g2_nand2_1 _13609_ (
    .A(_03380_),
    .B(_00269_),
    .Y(_03445_)
  );
  sg13g2_nand3_1 _13610_ (
    .A(_05247_),
    .B(_00884_),
    .C(_03445_),
    .Y(_03447_)
  );
  sg13g2_nor2_1 _13611_ (
    .A(_00112_),
    .B(_01580_),
    .Y(_03448_)
  );
  sg13g2_and2_1 _13612_ (
    .A(_03447_),
    .B(_03448_),
    .X(_03449_)
  );
  sg13g2_a21oi_1 _13613_ (
    .A1(_00083_),
    .A2(_01144_),
    .B1(addr_i_2_),
    .Y(_03450_)
  );
  sg13g2_o21ai_1 _13614_ (
    .A1(_03186_),
    .A2(_03450_),
    .B1(_01542_),
    .Y(_03451_)
  );
  sg13g2_nand2_1 _13615_ (
    .A(_00914_),
    .B(_02560_),
    .Y(_03452_)
  );
  sg13g2_nor2_1 _13616_ (
    .A(_01970_),
    .B(_03452_),
    .Y(_03453_)
  );
  sg13g2_nor4_1 _13617_ (
    .A(_04683_),
    .B(_00492_),
    .C(_00346_),
    .D(_03453_),
    .Y(_03454_)
  );
  sg13g2_buf_1 _13618_ (
    .A(_02423_),
    .X(_03455_)
  );
  sg13g2_nor4_1 _13619_ (
    .A(_01155_),
    .B(_01420_),
    .C(_03455_),
    .D(_02486_),
    .Y(_03456_)
  );
  sg13g2_nor2_1 _13620_ (
    .A(_05346_),
    .B(_00890_),
    .Y(_03458_)
  );
  sg13g2_o21ai_1 _13621_ (
    .A1(addr_i_4_),
    .A2(_00557_),
    .B1(_01432_),
    .Y(_03459_)
  );
  sg13g2_a21oi_1 _13622_ (
    .A1(_00371_),
    .A2(_01197_),
    .B1(addr_i_2_),
    .Y(_03460_)
  );
  sg13g2_a221oi_1 _13623_ (
    .A1(_00072_),
    .A2(_03458_),
    .B1(_03459_),
    .B2(addr_i_3_),
    .C1(_03460_),
    .Y(_03461_)
  );
  sg13g2_nor2_1 _13624_ (
    .A(_00351_),
    .B(_03461_),
    .Y(_03462_)
  );
  sg13g2_nor4_1 _13625_ (
    .A(addr_i_8_),
    .B(_03454_),
    .C(_03456_),
    .D(_03462_),
    .Y(_03463_)
  );
  sg13g2_a22oi_1 _13626_ (
    .A1(_03449_),
    .A2(_03451_),
    .B1(addr_i_9_),
    .B2(_03463_),
    .Y(_03464_)
  );
  sg13g2_nand2_1 _13627_ (
    .A(addr_i_8_),
    .B(addr_i_5_),
    .Y(_03465_)
  );
  sg13g2_nand2_1 _13628_ (
    .A(addr_i_7_),
    .B(_03465_),
    .Y(_03466_)
  );
  sg13g2_nand2_1 _13629_ (
    .A(addr_i_7_),
    .B(_05955_),
    .Y(_03467_)
  );
  sg13g2_nor2_1 _13630_ (
    .A(addr_i_3_),
    .B(_03467_),
    .Y(_03469_)
  );
  sg13g2_a22oi_1 _13631_ (
    .A1(addr_i_3_),
    .A2(_03466_),
    .B1(_03469_),
    .B2(_00243_),
    .Y(_03470_)
  );
  sg13g2_nor2_1 _13632_ (
    .A(_03464_),
    .B(_03470_),
    .Y(_03471_)
  );
  sg13g2_a21oi_1 _13633_ (
    .A1(_00703_),
    .A2(_04439_),
    .B1(_05833_),
    .Y(_03472_)
  );
  sg13g2_nand2b_1 _13634_ (
    .A_N(_03472_),
    .B(_00215_),
    .Y(_03473_)
  );
  sg13g2_o21ai_1 _13635_ (
    .A1(addr_i_10_),
    .A2(_03471_),
    .B1(_03473_),
    .Y(_03474_)
  );
  sg13g2_nor2_1 _13636_ (
    .A(_04837_),
    .B(_01402_),
    .Y(_03475_)
  );
  sg13g2_nor3_1 _13637_ (
    .A(addr_i_3_),
    .B(_00597_),
    .C(_00192_),
    .Y(_03476_)
  );
  sg13g2_a22oi_1 _13638_ (
    .A1(addr_i_3_),
    .A2(_03475_),
    .B1(_03476_),
    .B2(_06905_),
    .Y(_03477_)
  );
  sg13g2_nand2_1 _13639_ (
    .A(addr_i_6_),
    .B(_00008_),
    .Y(_03478_)
  );
  sg13g2_o21ai_1 _13640_ (
    .A1(addr_i_3_),
    .A2(_03478_),
    .B1(_00884_),
    .Y(_03480_)
  );
  sg13g2_o21ai_1 _13641_ (
    .A1(_03632_),
    .A2(_03523_),
    .B1(addr_i_3_),
    .Y(_03481_)
  );
  sg13g2_a21oi_1 _13642_ (
    .A1(_01694_),
    .A2(_03481_),
    .B1(_00122_),
    .Y(_03482_)
  );
  sg13g2_a21o_1 _13643_ (
    .A1(_01615_),
    .A2(_03480_),
    .B1(_03482_),
    .X(_03483_)
  );
  sg13g2_o21ai_1 _13644_ (
    .A1(_03477_),
    .A2(_03483_),
    .B1(_02604_),
    .Y(_03484_)
  );
  sg13g2_nand2_1 _13645_ (
    .A(addr_i_5_),
    .B(_01066_),
    .Y(_03485_)
  );
  sg13g2_nand3_1 _13646_ (
    .A(_01095_),
    .B(_01339_),
    .C(_03485_),
    .Y(_03486_)
  );
  sg13g2_a21oi_1 _13647_ (
    .A1(_02012_),
    .A2(_01168_),
    .B1(addr_i_3_),
    .Y(_03487_)
  );
  sg13g2_a21oi_1 _13648_ (
    .A1(_00582_),
    .A2(_00894_),
    .B1(_00083_),
    .Y(_03488_)
  );
  sg13g2_nor4_1 _13649_ (
    .A(_00128_),
    .B(_02535_),
    .C(_03487_),
    .D(_03488_),
    .Y(_03489_)
  );
  sg13g2_nand2_1 _13650_ (
    .A(_00355_),
    .B(_02954_),
    .Y(_03491_)
  );
  sg13g2_o21ai_1 _13651_ (
    .A1(_02443_),
    .A2(_01960_),
    .B1(_03491_),
    .Y(_03492_)
  );
  sg13g2_o21ai_1 _13652_ (
    .A1(_06276_),
    .A2(_00947_),
    .B1(addr_i_4_),
    .Y(_03493_)
  );
  sg13g2_nand2_1 _13653_ (
    .A(_05811_),
    .B(_00422_),
    .Y(_03494_)
  );
  sg13g2_a21oi_1 _13654_ (
    .A1(_03492_),
    .A2(_03493_),
    .B1(_03494_),
    .Y(_03495_)
  );
  sg13g2_a22oi_1 _13655_ (
    .A1(_03486_),
    .A2(_03489_),
    .B1(_03495_),
    .B2(addr_i_10_),
    .Y(_03496_)
  );
  sg13g2_buf_1 _13656_ (
    .A(_08941_),
    .X(_03497_)
  );
  sg13g2_a21oi_1 _13657_ (
    .A1(_00491_),
    .A2(_03497_),
    .B1(_01536_),
    .Y(_03498_)
  );
  sg13g2_o21ai_1 _13658_ (
    .A1(_00210_),
    .A2(_01243_),
    .B1(addr_i_4_),
    .Y(_03499_)
  );
  sg13g2_a21oi_1 _13659_ (
    .A1(_02799_),
    .A2(_03499_),
    .B1(_00006_),
    .Y(_03500_)
  );
  sg13g2_nand2_1 _13660_ (
    .A(addr_i_5_),
    .B(_07447_),
    .Y(_03502_)
  );
  sg13g2_a21oi_1 _13661_ (
    .A1(_03502_),
    .A2(_01463_),
    .B1(_00021_),
    .Y(_03503_)
  );
  sg13g2_a21oi_1 _13662_ (
    .A1(_01268_),
    .A2(_01389_),
    .B1(_00505_),
    .Y(_03504_)
  );
  sg13g2_nor4_1 _13663_ (
    .A(_06684_),
    .B(_03500_),
    .C(_03503_),
    .D(_03504_),
    .Y(_03505_)
  );
  sg13g2_o21ai_1 _13664_ (
    .A1(_00230_),
    .A2(_03498_),
    .B1(_03505_),
    .Y(_03506_)
  );
  sg13g2_a21oi_1 _13665_ (
    .A1(_00408_),
    .A2(_03324_),
    .B1(_02213_),
    .Y(_03507_)
  );
  sg13g2_a22oi_1 _13666_ (
    .A1(_00688_),
    .A2(_00641_),
    .B1(_03507_),
    .B2(addr_i_8_),
    .Y(_03508_)
  );
  sg13g2_nor2_1 _13667_ (
    .A(_02479_),
    .B(_07911_),
    .Y(_03509_)
  );
  sg13g2_o21ai_1 _13668_ (
    .A1(_07978_),
    .A2(_03509_),
    .B1(_00168_),
    .Y(_03510_)
  );
  sg13g2_nand3_1 _13669_ (
    .A(_02303_),
    .B(_03508_),
    .C(_03510_),
    .Y(_03511_)
  );
  sg13g2_nand3_1 _13670_ (
    .A(addr_i_9_),
    .B(_03506_),
    .C(_03511_),
    .Y(_03513_)
  );
  sg13g2_nand3_1 _13671_ (
    .A(_03484_),
    .B(_03496_),
    .C(_03513_),
    .Y(_03514_)
  );
  sg13g2_nand2_1 _13672_ (
    .A(addr_i_2_),
    .B(_01037_),
    .Y(_03515_)
  );
  sg13g2_or3_1 _13673_ (
    .A(addr_i_2_),
    .B(_00119_),
    .C(_00204_),
    .X(_03516_)
  );
  sg13g2_o21ai_1 _13674_ (
    .A1(_02937_),
    .A2(_03515_),
    .B1(_03516_),
    .Y(_03517_)
  );
  sg13g2_o21ai_1 _13675_ (
    .A1(_02343_),
    .A2(_02395_),
    .B1(_00938_),
    .Y(_03518_)
  );
  sg13g2_nand2_1 _13676_ (
    .A(_05943_),
    .B(_03676_),
    .Y(_03519_)
  );
  sg13g2_nand2_1 _13677_ (
    .A(addr_i_7_),
    .B(_03519_),
    .Y(_03520_)
  );
  sg13g2_o21ai_1 _13678_ (
    .A1(_05424_),
    .A2(_07193_),
    .B1(addr_i_3_),
    .Y(_03521_)
  );
  sg13g2_a21oi_1 _13679_ (
    .A1(_00131_),
    .A2(_03521_),
    .B1(addr_i_4_),
    .Y(_03522_)
  );
  sg13g2_a22oi_1 _13680_ (
    .A1(addr_i_4_),
    .A2(_03518_),
    .B1(_03520_),
    .B2(_03522_),
    .Y(_03524_)
  );
  sg13g2_a21oi_1 _13681_ (
    .A1(_01615_),
    .A2(_03517_),
    .B1(_03524_),
    .Y(_03525_)
  );
  sg13g2_nand2_1 _13682_ (
    .A(_01310_),
    .B(_01354_),
    .Y(_03526_)
  );
  sg13g2_o21ai_1 _13683_ (
    .A1(_06176_),
    .A2(_00205_),
    .B1(addr_i_3_),
    .Y(_03527_)
  );
  sg13g2_o21ai_1 _13684_ (
    .A1(addr_i_6_),
    .A2(_09484_),
    .B1(_03527_),
    .Y(_03528_)
  );
  sg13g2_nand2_1 _13685_ (
    .A(_01589_),
    .B(_07922_),
    .Y(_03529_)
  );
  sg13g2_a21oi_1 _13686_ (
    .A1(_05036_),
    .A2(_00571_),
    .B1(addr_i_3_),
    .Y(_03530_)
  );
  sg13g2_a22oi_1 _13687_ (
    .A1(_03245_),
    .A2(_08033_),
    .B1(_03529_),
    .B2(_03530_),
    .Y(_03531_)
  );
  sg13g2_o21ai_1 _13688_ (
    .A1(_08598_),
    .A2(_01144_),
    .B1(_03531_),
    .Y(_03532_)
  );
  sg13g2_o21ai_1 _13689_ (
    .A1(_03526_),
    .A2(_03528_),
    .B1(_03532_),
    .Y(_03533_)
  );
  sg13g2_a22oi_1 _13690_ (
    .A1(_00782_),
    .A2(_03525_),
    .B1(_03533_),
    .B2(_02700_),
    .Y(_03535_)
  );
  sg13g2_a21o_1 _13691_ (
    .A1(addr_i_2_),
    .A2(_00194_),
    .B1(_02388_),
    .X(_03536_)
  );
  sg13g2_nor3_1 _13692_ (
    .A(_07491_),
    .B(addr_i_5_),
    .C(_01680_),
    .Y(_03537_)
  );
  sg13g2_a21oi_1 _13693_ (
    .A1(_08221_),
    .A2(_00618_),
    .B1(_03765_),
    .Y(_03538_)
  );
  sg13g2_or2_1 _13694_ (
    .A(_03537_),
    .B(_03538_),
    .X(_03539_)
  );
  sg13g2_buf_1 _13695_ (
    .A(_00245_),
    .X(_03540_)
  );
  sg13g2_o21ai_1 _13696_ (
    .A1(addr_i_4_),
    .A2(_01507_),
    .B1(_03540_),
    .Y(_03541_)
  );
  sg13g2_nand2_1 _13697_ (
    .A(addr_i_3_),
    .B(_01740_),
    .Y(_03542_)
  );
  sg13g2_a221oi_1 _13698_ (
    .A1(addr_i_4_),
    .A2(_03539_),
    .B1(_03541_),
    .B2(_00534_),
    .C1(_03542_),
    .Y(_03543_)
  );
  sg13g2_a22oi_1 _13699_ (
    .A1(_00047_),
    .A2(_03536_),
    .B1(_03543_),
    .B2(addr_i_8_),
    .Y(_03544_)
  );
  sg13g2_nand2_1 _13700_ (
    .A(_00477_),
    .B(_01715_),
    .Y(_03546_)
  );
  sg13g2_a22oi_1 _13701_ (
    .A1(addr_i_3_),
    .A2(_03546_),
    .B1(_03720_),
    .B2(_00491_),
    .Y(_03547_)
  );
  sg13g2_nor3_1 _13702_ (
    .A(_05932_),
    .B(_00009_),
    .C(_01777_),
    .Y(_03548_)
  );
  sg13g2_a22oi_1 _13703_ (
    .A1(_00319_),
    .A2(_00702_),
    .B1(_01494_),
    .B2(_02598_),
    .Y(_03549_)
  );
  sg13g2_o21ai_1 _13704_ (
    .A1(addr_i_2_),
    .A2(_03548_),
    .B1(_03549_),
    .Y(_03550_)
  );
  sg13g2_o21ai_1 _13705_ (
    .A1(_03227_),
    .A2(_03547_),
    .B1(_03550_),
    .Y(_03551_)
  );
  sg13g2_nor3_1 _13706_ (
    .A(addr_i_9_),
    .B(_03544_),
    .C(_03551_),
    .Y(_03552_)
  );
  sg13g2_o21ai_1 _13707_ (
    .A1(_03535_),
    .A2(_03552_),
    .B1(addr_i_10_),
    .Y(_03553_)
  );
  sg13g2_and2_1 _13708_ (
    .A(_03514_),
    .B(_03553_),
    .X(_03554_)
  );
  sg13g2_mux4_1 _13709_ (
    .A0(_03356_),
    .A1(_03444_),
    .A2(_03474_),
    .A3(_03554_),
    .S0(_03051_),
    .S1(addr_i_12_),
    .X(data_o_18_)
  );
  sg13g2_nor2_1 _13710_ (
    .A(addr_i_5_),
    .B(_04218_),
    .Y(_03556_)
  );
  sg13g2_nand2_1 _13711_ (
    .A(_00304_),
    .B(_03556_),
    .Y(_03557_)
  );
  sg13g2_o21ai_1 _13712_ (
    .A1(_00105_),
    .A2(_02289_),
    .B1(_03557_),
    .Y(_03558_)
  );
  sg13g2_nand2_1 _13713_ (
    .A(_00483_),
    .B(_03110_),
    .Y(_03559_)
  );
  sg13g2_a22oi_1 _13714_ (
    .A1(_09260_),
    .A2(_03559_),
    .B1(addr_i_4_),
    .B2(_03238_),
    .Y(_03560_)
  );
  sg13g2_a22oi_1 _13715_ (
    .A1(_00440_),
    .A2(_03558_),
    .B1(_03560_),
    .B2(_00397_),
    .Y(_03561_)
  );
  sg13g2_nor2_1 _13716_ (
    .A(_04793_),
    .B(_01899_),
    .Y(_03562_)
  );
  sg13g2_a21o_1 _13717_ (
    .A1(_00542_),
    .A2(_00842_),
    .B1(_03562_),
    .X(_03563_)
  );
  sg13g2_o21ai_1 _13718_ (
    .A1(_02042_),
    .A2(_01091_),
    .B1(addr_i_3_),
    .Y(_03564_)
  );
  sg13g2_nor2_1 _13719_ (
    .A(_00327_),
    .B(_01636_),
    .Y(_03565_)
  );
  sg13g2_o21ai_1 _13720_ (
    .A1(_02265_),
    .A2(_03565_),
    .B1(_05877_),
    .Y(_03567_)
  );
  sg13g2_a21oi_1 _13721_ (
    .A1(_03564_),
    .A2(_03567_),
    .B1(_01391_),
    .Y(_03568_)
  );
  sg13g2_a21oi_1 _13722_ (
    .A1(_00277_),
    .A2(_03563_),
    .B1(_03568_),
    .Y(_03569_)
  );
  sg13g2_nand2_1 _13723_ (
    .A(addr_i_3_),
    .B(_01033_),
    .Y(_03570_)
  );
  sg13g2_a22oi_1 _13724_ (
    .A1(_00467_),
    .A2(_03570_),
    .B1(_00747_),
    .B2(_08487_),
    .Y(_03571_)
  );
  sg13g2_buf_1 _13725_ (
    .A(_02153_),
    .X(_03572_)
  );
  sg13g2_a21oi_1 _13726_ (
    .A1(addr_i_3_),
    .A2(_02214_),
    .B1(_02639_),
    .Y(_03573_)
  );
  sg13g2_nor2_1 _13727_ (
    .A(addr_i_2_),
    .B(_03573_),
    .Y(_03574_)
  );
  sg13g2_buf_1 _13728_ (
    .A(_04715_),
    .X(_03575_)
  );
  sg13g2_xnor2_1 _13729_ (
    .A(_04981_),
    .B(_00702_),
    .Y(_03576_)
  );
  sg13g2_a21oi_1 _13730_ (
    .A1(_03575_),
    .A2(_03576_),
    .B1(_00070_),
    .Y(_03578_)
  );
  sg13g2_a22oi_1 _13731_ (
    .A1(_01240_),
    .A2(_03572_),
    .B1(_03574_),
    .B2(_03578_),
    .Y(_03579_)
  );
  sg13g2_nor2_1 _13732_ (
    .A(addr_i_8_),
    .B(_03579_),
    .Y(_03580_)
  );
  sg13g2_nand2_1 _13733_ (
    .A(_02598_),
    .B(_00960_),
    .Y(_03581_)
  );
  sg13g2_o21ai_1 _13734_ (
    .A1(_01024_),
    .A2(_07967_),
    .B1(_05711_),
    .Y(_03582_)
  );
  sg13g2_a21o_1 _13735_ (
    .A1(_00414_),
    .A2(_03582_),
    .B1(addr_i_5_),
    .X(_03583_)
  );
  sg13g2_a21oi_1 _13736_ (
    .A1(_03581_),
    .A2(_03583_),
    .B1(_01391_),
    .Y(_03584_)
  );
  sg13g2_nor4_1 _13737_ (
    .A(addr_i_9_),
    .B(_03571_),
    .C(_03580_),
    .D(_03584_),
    .Y(_03585_)
  );
  sg13g2_a21oi_1 _13738_ (
    .A1(_03561_),
    .A2(_03569_),
    .B1(_03585_),
    .Y(_03586_)
  );
  sg13g2_nor2_1 _13739_ (
    .A(_01065_),
    .B(_00079_),
    .Y(_03587_)
  );
  sg13g2_nor2_1 _13740_ (
    .A(_07602_),
    .B(_02031_),
    .Y(_03589_)
  );
  sg13g2_o21ai_1 _13741_ (
    .A1(_03587_),
    .A2(_03589_),
    .B1(addr_i_3_),
    .Y(_03590_)
  );
  sg13g2_o21ai_1 _13742_ (
    .A1(_02349_),
    .A2(_02578_),
    .B1(_03590_),
    .Y(_03591_)
  );
  sg13g2_nor2_1 _13743_ (
    .A(_00172_),
    .B(_02368_),
    .Y(_03592_)
  );
  sg13g2_a22oi_1 _13744_ (
    .A1(_02832_),
    .A2(_01230_),
    .B1(_03203_),
    .B2(_00151_),
    .Y(_03593_)
  );
  sg13g2_o21ai_1 _13745_ (
    .A1(_01660_),
    .A2(_04837_),
    .B1(addr_i_3_),
    .Y(_03594_)
  );
  sg13g2_a21oi_1 _13746_ (
    .A1(_01336_),
    .A2(_00118_),
    .B1(_00399_),
    .Y(_03595_)
  );
  sg13g2_a21oi_1 _13747_ (
    .A1(_03594_),
    .A2(_03595_),
    .B1(_02963_),
    .Y(_03596_)
  );
  sg13g2_a22oi_1 _13748_ (
    .A1(_03591_),
    .A2(_03592_),
    .B1(_03593_),
    .B2(_03596_),
    .Y(_03597_)
  );
  sg13g2_nand2_1 _13749_ (
    .A(_00818_),
    .B(_01923_),
    .Y(_03598_)
  );
  sg13g2_nand3_1 _13750_ (
    .A(addr_i_8_),
    .B(_07824_),
    .C(_00688_),
    .Y(_03600_)
  );
  sg13g2_nor2_1 _13751_ (
    .A(_00064_),
    .B(_05955_),
    .Y(_03601_)
  );
  sg13g2_o21ai_1 _13752_ (
    .A1(_01107_),
    .A2(_03601_),
    .B1(addr_i_3_),
    .Y(_03602_)
  );
  sg13g2_nand3_1 _13753_ (
    .A(_03598_),
    .B(_03600_),
    .C(_03602_),
    .Y(_03603_)
  );
  sg13g2_o21ai_1 _13754_ (
    .A1(_03632_),
    .A2(_00177_),
    .B1(addr_i_3_),
    .Y(_03604_)
  );
  sg13g2_a21oi_1 _13755_ (
    .A1(_01425_),
    .A2(_03604_),
    .B1(addr_i_8_),
    .Y(_03605_)
  );
  sg13g2_a21oi_1 _13756_ (
    .A1(addr_i_8_),
    .A2(_08598_),
    .B1(_01420_),
    .Y(_03606_)
  );
  sg13g2_nor2b_1 _13757_ (
    .A(addr_i_3_),
    .B_N(addr_i_8_),
    .Y(_03607_)
  );
  sg13g2_a21oi_1 _13758_ (
    .A1(_02055_),
    .A2(_03607_),
    .B1(_01615_),
    .Y(_03608_)
  );
  sg13g2_o21ai_1 _13759_ (
    .A1(_00943_),
    .A2(_03606_),
    .B1(_03608_),
    .Y(_03609_)
  );
  sg13g2_a22oi_1 _13760_ (
    .A1(addr_i_6_),
    .A2(_03603_),
    .B1(_03605_),
    .B2(_03609_),
    .Y(_03611_)
  );
  sg13g2_a21oi_1 _13761_ (
    .A1(addr_i_3_),
    .A2(_06441_),
    .B1(_06320_),
    .Y(_03612_)
  );
  sg13g2_nand3_1 _13762_ (
    .A(_09491_),
    .B(_02815_),
    .C(_03465_),
    .Y(_03613_)
  );
  sg13g2_o21ai_1 _13763_ (
    .A1(addr_i_6_),
    .A2(_03612_),
    .B1(_03613_),
    .Y(_03614_)
  );
  sg13g2_nor3_1 _13764_ (
    .A(addr_i_8_),
    .B(_00128_),
    .C(_07558_),
    .Y(_03615_)
  );
  sg13g2_a22oi_1 _13765_ (
    .A1(addr_i_2_),
    .A2(_03614_),
    .B1(_03615_),
    .B2(addr_i_4_),
    .Y(_03616_)
  );
  sg13g2_buf_1 _13766_ (
    .A(_01548_),
    .X(_03617_)
  );
  sg13g2_nor3_1 _13767_ (
    .A(_08785_),
    .B(addr_i_5_),
    .C(_01917_),
    .Y(_03618_)
  );
  sg13g2_nor2_1 _13768_ (
    .A(_01548_),
    .B(_03743_),
    .Y(_03619_)
  );
  sg13g2_or2_1 _13769_ (
    .A(_03618_),
    .B(_03619_),
    .X(_03620_)
  );
  sg13g2_a221oi_1 _13770_ (
    .A1(_03617_),
    .A2(_02170_),
    .B1(_03620_),
    .B2(addr_i_2_),
    .C1(_01794_),
    .Y(_03622_)
  );
  sg13g2_a21oi_1 _13771_ (
    .A1(_01480_),
    .A2(_01920_),
    .B1(addr_i_7_),
    .Y(_03623_)
  );
  sg13g2_o21ai_1 _13772_ (
    .A1(_03616_),
    .A2(_03622_),
    .B1(_03623_),
    .Y(_03624_)
  );
  sg13g2_nand3b_1 _13773_ (
    .A_N(_03611_),
    .B(_03624_),
    .C(addr_i_9_),
    .Y(_03625_)
  );
  sg13g2_a21oi_1 _13774_ (
    .A1(_03597_),
    .A2(_03625_),
    .B1(addr_i_10_),
    .Y(_03626_)
  );
  sg13g2_a22oi_1 _13775_ (
    .A1(addr_i_10_),
    .A2(_03586_),
    .B1(_03626_),
    .B2(addr_i_11_),
    .Y(_03627_)
  );
  sg13g2_a21oi_1 _13776_ (
    .A1(_00070_),
    .A2(_02254_),
    .B1(_00185_),
    .Y(_03628_)
  );
  sg13g2_a21oi_1 _13777_ (
    .A1(_01508_),
    .A2(_01765_),
    .B1(_03628_),
    .Y(_03629_)
  );
  sg13g2_o21ai_1 _13778_ (
    .A1(_01277_),
    .A2(_05645_),
    .B1(addr_i_4_),
    .Y(_03630_)
  );
  sg13g2_nor2_1 _13779_ (
    .A(_03798_),
    .B(_00664_),
    .Y(_03631_)
  );
  sg13g2_o21ai_1 _13780_ (
    .A1(_03643_),
    .A2(_03631_),
    .B1(addr_i_2_),
    .Y(_03633_)
  );
  sg13g2_a21oi_1 _13781_ (
    .A1(_03630_),
    .A2(_03633_),
    .B1(addr_i_3_),
    .Y(_03634_)
  );
  sg13g2_a21oi_1 _13782_ (
    .A1(_00500_),
    .A2(_03572_),
    .B1(_03634_),
    .Y(_03635_)
  );
  sg13g2_o21ai_1 _13783_ (
    .A1(_00048_),
    .A2(_03629_),
    .B1(_03635_),
    .Y(_03636_)
  );
  sg13g2_a21oi_1 _13784_ (
    .A1(addr_i_2_),
    .A2(_04616_),
    .B1(_00231_),
    .Y(_03637_)
  );
  sg13g2_a21oi_1 _13785_ (
    .A1(_03091_),
    .A2(_03273_),
    .B1(addr_i_6_),
    .Y(_03638_)
  );
  sg13g2_a221oi_1 _13786_ (
    .A1(_00022_),
    .A2(_01227_),
    .B1(_03637_),
    .B2(_01240_),
    .C1(_03638_),
    .Y(_03639_)
  );
  sg13g2_a21oi_1 _13787_ (
    .A1(addr_i_3_),
    .A2(_00282_),
    .B1(_08299_),
    .Y(_03640_)
  );
  sg13g2_o21ai_1 _13788_ (
    .A1(addr_i_4_),
    .A2(_03640_),
    .B1(_00739_),
    .Y(_03641_)
  );
  sg13g2_nor2_1 _13789_ (
    .A(addr_i_7_),
    .B(_03641_),
    .Y(_03642_)
  );
  sg13g2_a22oi_1 _13790_ (
    .A1(addr_i_7_),
    .A2(_03639_),
    .B1(_03642_),
    .B2(addr_i_8_),
    .Y(_03644_)
  );
  sg13g2_a22oi_1 _13791_ (
    .A1(addr_i_8_),
    .A2(_03636_),
    .B1(_03644_),
    .B2(addr_i_9_),
    .Y(_03645_)
  );
  sg13g2_o21ai_1 _13792_ (
    .A1(_07757_),
    .A2(_00205_),
    .B1(addr_i_3_),
    .Y(_03646_)
  );
  sg13g2_a21oi_1 _13793_ (
    .A1(_00368_),
    .A2(_03646_),
    .B1(addr_i_2_),
    .Y(_03647_)
  );
  sg13g2_nor2_1 _13794_ (
    .A(_09038_),
    .B(_00078_),
    .Y(_03648_)
  );
  sg13g2_a22oi_1 _13795_ (
    .A1(_08785_),
    .A2(_09215_),
    .B1(_03648_),
    .B2(_01107_),
    .Y(_03649_)
  );
  sg13g2_o21ai_1 _13796_ (
    .A1(addr_i_6_),
    .A2(_03649_),
    .B1(addr_i_7_),
    .Y(_03650_)
  );
  sg13g2_or2_1 _13797_ (
    .A(_03647_),
    .B(_03650_),
    .X(_03651_)
  );
  sg13g2_buf_1 _13798_ (
    .A(_00354_),
    .X(_03652_)
  );
  sg13g2_o21ai_1 _13799_ (
    .A1(addr_i_3_),
    .A2(_01789_),
    .B1(_01527_),
    .Y(_03653_)
  );
  sg13g2_a22oi_1 _13800_ (
    .A1(_03652_),
    .A2(_03653_),
    .B1(_03562_),
    .B2(addr_i_7_),
    .Y(_03655_)
  );
  sg13g2_nor2_1 _13801_ (
    .A(addr_i_8_),
    .B(_03655_),
    .Y(_03656_)
  );
  sg13g2_o21ai_1 _13802_ (
    .A1(addr_i_6_),
    .A2(_04097_),
    .B1(_01353_),
    .Y(_03657_)
  );
  sg13g2_nor2_1 _13803_ (
    .A(_00522_),
    .B(_01789_),
    .Y(_03658_)
  );
  sg13g2_a21oi_1 _13804_ (
    .A1(addr_i_4_),
    .A2(_03657_),
    .B1(_03658_),
    .Y(_03659_)
  );
  sg13g2_nand2_1 _13805_ (
    .A(_00593_),
    .B(_07757_),
    .Y(_03660_)
  );
  sg13g2_o21ai_1 _13806_ (
    .A1(_00046_),
    .A2(_03258_),
    .B1(_03660_),
    .Y(_03661_)
  );
  sg13g2_nand2_1 _13807_ (
    .A(_08930_),
    .B(_01197_),
    .Y(_03662_)
  );
  sg13g2_nor2_1 _13808_ (
    .A(_02472_),
    .B(_03662_),
    .Y(_03663_)
  );
  sg13g2_a22oi_1 _13809_ (
    .A1(addr_i_2_),
    .A2(_03661_),
    .B1(_03663_),
    .B2(addr_i_7_),
    .Y(_03664_)
  );
  sg13g2_a22oi_1 _13810_ (
    .A1(addr_i_7_),
    .A2(_03659_),
    .B1(_03664_),
    .B2(_01043_),
    .Y(_03666_)
  );
  sg13g2_a22oi_1 _13811_ (
    .A1(_03651_),
    .A2(_03656_),
    .B1(_01351_),
    .B2(_03666_),
    .Y(_03667_)
  );
  sg13g2_or2_1 _13812_ (
    .A(addr_i_10_),
    .B(_03667_),
    .X(_03668_)
  );
  sg13g2_nand2_1 _13813_ (
    .A(_08785_),
    .B(_00578_),
    .Y(_03669_)
  );
  sg13g2_nand3_1 _13814_ (
    .A(addr_i_4_),
    .B(_00736_),
    .C(_00938_),
    .Y(_03670_)
  );
  sg13g2_nor2_1 _13815_ (
    .A(_00479_),
    .B(_04683_),
    .Y(_03671_)
  );
  sg13g2_nand2_1 _13816_ (
    .A(_03670_),
    .B(_03671_),
    .Y(_03672_)
  );
  sg13g2_a21oi_1 _13817_ (
    .A1(_03669_),
    .A2(_03672_),
    .B1(_03227_),
    .Y(_03673_)
  );
  sg13g2_a21oi_1 _13818_ (
    .A1(_05546_),
    .A2(_02799_),
    .B1(addr_i_3_),
    .Y(_03674_)
  );
  sg13g2_o21ai_1 _13819_ (
    .A1(_00850_),
    .A2(_03674_),
    .B1(addr_i_6_),
    .Y(_03675_)
  );
  sg13g2_o21ai_1 _13820_ (
    .A1(_01120_),
    .A2(_00993_),
    .B1(_01432_),
    .Y(_03677_)
  );
  sg13g2_a21oi_1 _13821_ (
    .A1(addr_i_3_),
    .A2(_03677_),
    .B1(_01402_),
    .Y(_03678_)
  );
  sg13g2_a21oi_1 _13822_ (
    .A1(_03675_),
    .A2(_03678_),
    .B1(_08674_),
    .Y(_03679_)
  );
  sg13g2_nand2_1 _13823_ (
    .A(_01589_),
    .B(_00852_),
    .Y(_03680_)
  );
  sg13g2_o21ai_1 _13824_ (
    .A1(_09172_),
    .A2(_03680_),
    .B1(addr_i_5_),
    .Y(_03681_)
  );
  sg13g2_a21o_1 _13825_ (
    .A1(addr_i_3_),
    .A2(_03170_),
    .B1(_01093_),
    .X(_03682_)
  );
  sg13g2_a22oi_1 _13826_ (
    .A1(addr_i_4_),
    .A2(_03682_),
    .B1(_00587_),
    .B2(addr_i_7_),
    .Y(_03683_)
  );
  sg13g2_nand2_1 _13827_ (
    .A(_00137_),
    .B(_01912_),
    .Y(_03684_)
  );
  sg13g2_a21oi_1 _13828_ (
    .A1(_04063_),
    .A2(_01197_),
    .B1(addr_i_6_),
    .Y(_03685_)
  );
  sg13g2_a22oi_1 _13829_ (
    .A1(_02990_),
    .A2(_03684_),
    .B1(_03685_),
    .B2(_02424_),
    .Y(_03686_)
  );
  sg13g2_a221oi_1 _13830_ (
    .A1(_03681_),
    .A2(_03683_),
    .B1(_03686_),
    .B2(addr_i_7_),
    .C1(addr_i_8_),
    .Y(_03688_)
  );
  sg13g2_or3_1 _13831_ (
    .A(_03673_),
    .B(_03679_),
    .C(_03688_),
    .X(_03689_)
  );
  sg13g2_buf_1 _13832_ (
    .A(_00099_),
    .X(_03690_)
  );
  sg13g2_nor3_1 _13833_ (
    .A(addr_i_3_),
    .B(_05280_),
    .C(_03690_),
    .Y(_03691_)
  );
  sg13g2_nor2_1 _13834_ (
    .A(addr_i_4_),
    .B(_01228_),
    .Y(_03692_)
  );
  sg13g2_a22oi_1 _13835_ (
    .A1(_01065_),
    .A2(_00960_),
    .B1(_03692_),
    .B2(addr_i_2_),
    .Y(_03693_)
  );
  sg13g2_or4_1 _13836_ (
    .A(addr_i_6_),
    .B(_02327_),
    .C(_03691_),
    .D(_03693_),
    .X(_03694_)
  );
  sg13g2_nor2_1 _13837_ (
    .A(addr_i_4_),
    .B(_01652_),
    .Y(_03695_)
  );
  sg13g2_o21ai_1 _13838_ (
    .A1(_02734_),
    .A2(_03695_),
    .B1(_01508_),
    .Y(_03696_)
  );
  sg13g2_a21oi_1 _13839_ (
    .A1(addr_i_3_),
    .A2(_04429_),
    .B1(_03380_),
    .Y(_03697_)
  );
  sg13g2_nor2_1 _13840_ (
    .A(_00293_),
    .B(_03697_),
    .Y(_03699_)
  );
  sg13g2_o21ai_1 _13841_ (
    .A1(_01192_),
    .A2(_03699_),
    .B1(addr_i_6_),
    .Y(_03700_)
  );
  sg13g2_nand2_1 _13842_ (
    .A(_01881_),
    .B(_01972_),
    .Y(_03701_)
  );
  sg13g2_a21o_1 _13843_ (
    .A1(_03700_),
    .A2(_03701_),
    .B1(addr_i_2_),
    .X(_03702_)
  );
  sg13g2_nand4_1 _13844_ (
    .A(addr_i_8_),
    .B(_03694_),
    .C(_03696_),
    .D(_03702_),
    .Y(_03703_)
  );
  sg13g2_a21oi_1 _13845_ (
    .A1(_00032_),
    .A2(_00404_),
    .B1(_00034_),
    .Y(_03704_)
  );
  sg13g2_a22oi_1 _13846_ (
    .A1(addr_i_4_),
    .A2(_01338_),
    .B1(_03704_),
    .B2(_00569_),
    .Y(_03705_)
  );
  sg13g2_a21oi_1 _13847_ (
    .A1(addr_i_3_),
    .A2(_00965_),
    .B1(_03033_),
    .Y(_03706_)
  );
  sg13g2_nand2_1 _13848_ (
    .A(_09050_),
    .B(_01243_),
    .Y(_03707_)
  );
  sg13g2_o21ai_1 _13849_ (
    .A1(_06607_),
    .A2(_03706_),
    .B1(_03707_),
    .Y(_03708_)
  );
  sg13g2_nand2_1 _13850_ (
    .A(_03380_),
    .B(_00454_),
    .Y(_03710_)
  );
  sg13g2_a21oi_1 _13851_ (
    .A1(_00055_),
    .A2(_03710_),
    .B1(addr_i_6_),
    .Y(_03711_)
  );
  sg13g2_a22oi_1 _13852_ (
    .A1(addr_i_2_),
    .A2(_03708_),
    .B1(_03711_),
    .B2(addr_i_8_),
    .Y(_03712_)
  );
  sg13g2_o21ai_1 _13853_ (
    .A1(addr_i_2_),
    .A2(_03705_),
    .B1(_03712_),
    .Y(_03713_)
  );
  sg13g2_and2_1 _13854_ (
    .A(_05203_),
    .B(_03713_),
    .X(_03714_)
  );
  sg13g2_a221oi_1 _13855_ (
    .A1(_01174_),
    .A2(_03689_),
    .B1(_03703_),
    .B2(_03714_),
    .C1(_03040_),
    .Y(_03715_)
  );
  sg13g2_o21ai_1 _13856_ (
    .A1(_03645_),
    .A2(_03668_),
    .B1(_03715_),
    .Y(_03716_)
  );
  sg13g2_nand2_1 _13857_ (
    .A(_02251_),
    .B(_03716_),
    .Y(_03717_)
  );
  sg13g2_a22oi_1 _13858_ (
    .A1(_00223_),
    .A2(_00301_),
    .B1(_00026_),
    .B2(_01559_),
    .Y(_03718_)
  );
  sg13g2_o21ai_1 _13859_ (
    .A1(_01199_),
    .A2(_00719_),
    .B1(_00656_),
    .Y(_03719_)
  );
  sg13g2_nand2_1 _13860_ (
    .A(_01658_),
    .B(_00413_),
    .Y(_03721_)
  );
  sg13g2_a22oi_1 _13861_ (
    .A1(_00463_),
    .A2(_03721_),
    .B1(_01319_),
    .B2(addr_i_5_),
    .Y(_03722_)
  );
  sg13g2_nand2_1 _13862_ (
    .A(_01965_),
    .B(_00618_),
    .Y(_03723_)
  );
  sg13g2_a22oi_1 _13863_ (
    .A1(addr_i_3_),
    .A2(_03723_),
    .B1(_02983_),
    .B2(_02874_),
    .Y(_03724_)
  );
  sg13g2_o21ai_1 _13864_ (
    .A1(_03722_),
    .A2(_03724_),
    .B1(addr_i_4_),
    .Y(_03725_)
  );
  sg13g2_o21ai_1 _13865_ (
    .A1(addr_i_4_),
    .A2(_03719_),
    .B1(_03725_),
    .Y(_03726_)
  );
  sg13g2_o21ai_1 _13866_ (
    .A1(_04296_),
    .A2(_01103_),
    .B1(_01004_),
    .Y(_03727_)
  );
  sg13g2_nand2_1 _13867_ (
    .A(_00112_),
    .B(_00633_),
    .Y(_03728_)
  );
  sg13g2_o21ai_1 _13868_ (
    .A1(_06972_),
    .A2(_08564_),
    .B1(_02799_),
    .Y(_03729_)
  );
  sg13g2_nor2_1 _13869_ (
    .A(_02471_),
    .B(_00543_),
    .Y(_03730_)
  );
  sg13g2_a21oi_1 _13870_ (
    .A1(addr_i_3_),
    .A2(_03729_),
    .B1(_03730_),
    .Y(_03733_)
  );
  sg13g2_nor2_1 _13871_ (
    .A(addr_i_6_),
    .B(_03733_),
    .Y(_03734_)
  );
  sg13g2_a22oi_1 _13872_ (
    .A1(_02277_),
    .A2(_03727_),
    .B1(_03728_),
    .B2(_03734_),
    .Y(_03735_)
  );
  sg13g2_a22oi_1 _13873_ (
    .A1(_03718_),
    .A2(_03726_),
    .B1(_03735_),
    .B2(addr_i_9_),
    .Y(_03736_)
  );
  sg13g2_nand2_1 _13874_ (
    .A(_07326_),
    .B(_03139_),
    .Y(_03737_)
  );
  sg13g2_o21ai_1 _13875_ (
    .A1(_04373_),
    .A2(_00745_),
    .B1(_03737_),
    .Y(_03738_)
  );
  sg13g2_o21ai_1 _13876_ (
    .A1(_06099_),
    .A2(_06563_),
    .B1(addr_i_4_),
    .Y(_03739_)
  );
  sg13g2_nand3_1 _13877_ (
    .A(addr_i_3_),
    .B(_01354_),
    .C(_03739_),
    .Y(_03740_)
  );
  sg13g2_o21ai_1 _13878_ (
    .A1(addr_i_3_),
    .A2(_03738_),
    .B1(_03740_),
    .Y(_03741_)
  );
  sg13g2_nor2_1 _13879_ (
    .A(_01757_),
    .B(_08453_),
    .Y(_03742_)
  );
  sg13g2_nor4_1 _13880_ (
    .A(_03186_),
    .B(_00866_),
    .C(_03562_),
    .D(_03742_),
    .Y(_03744_)
  );
  sg13g2_nand2_1 _13881_ (
    .A(_04151_),
    .B(_08288_),
    .Y(_03745_)
  );
  sg13g2_nand2_1 _13882_ (
    .A(_03665_),
    .B(_00158_),
    .Y(_03746_)
  );
  sg13g2_nand4_1 _13883_ (
    .A(_03391_),
    .B(_03744_),
    .C(_03745_),
    .D(_03746_),
    .Y(_03747_)
  );
  sg13g2_a22oi_1 _13884_ (
    .A1(_00380_),
    .A2(_02031_),
    .B1(_00210_),
    .B2(_00435_),
    .Y(_03748_)
  );
  sg13g2_a22oi_1 _13885_ (
    .A1(_06143_),
    .A2(_00030_),
    .B1(_00316_),
    .B2(_01888_),
    .Y(_03749_)
  );
  sg13g2_or2_1 _13886_ (
    .A(_03748_),
    .B(_03749_),
    .X(_03750_)
  );
  sg13g2_a22oi_1 _13887_ (
    .A1(addr_i_7_),
    .A2(_03747_),
    .B1(_03750_),
    .B2(addr_i_8_),
    .Y(_03751_)
  );
  sg13g2_nand3_1 _13888_ (
    .A(_01310_),
    .B(_02810_),
    .C(_03557_),
    .Y(_03752_)
  );
  sg13g2_nand2_1 _13889_ (
    .A(addr_i_3_),
    .B(_02181_),
    .Y(_03753_)
  );
  sg13g2_o21ai_1 _13890_ (
    .A1(_01103_),
    .A2(_01539_),
    .B1(_03753_),
    .Y(_03755_)
  );
  sg13g2_o21ai_1 _13891_ (
    .A1(_03752_),
    .A2(_03755_),
    .B1(addr_i_9_),
    .Y(_03756_)
  );
  sg13g2_a22oi_1 _13892_ (
    .A1(_00708_),
    .A2(_03741_),
    .B1(_03751_),
    .B2(_03756_),
    .Y(_03757_)
  );
  sg13g2_or3_1 _13893_ (
    .A(addr_i_10_),
    .B(_03736_),
    .C(_03757_),
    .X(_03758_)
  );
  sg13g2_nor2_1 _13894_ (
    .A(_02196_),
    .B(_01757_),
    .Y(_03759_)
  );
  sg13g2_a22oi_1 _13895_ (
    .A1(_00783_),
    .A2(_00666_),
    .B1(_03759_),
    .B2(addr_i_4_),
    .Y(_03760_)
  );
  sg13g2_nand2_1 _13896_ (
    .A(addr_i_6_),
    .B(_00495_),
    .Y(_03761_)
  );
  sg13g2_nor2_1 _13897_ (
    .A(addr_i_3_),
    .B(_03761_),
    .Y(_03762_)
  );
  sg13g2_a22oi_1 _13898_ (
    .A1(addr_i_3_),
    .A2(_09448_),
    .B1(_03762_),
    .B2(_09271_),
    .Y(_03763_)
  );
  sg13g2_nor3_1 _13899_ (
    .A(_08830_),
    .B(_03760_),
    .C(_03763_),
    .Y(_03764_)
  );
  sg13g2_o21ai_1 _13900_ (
    .A1(addr_i_2_),
    .A2(_00539_),
    .B1(_06485_),
    .Y(_03766_)
  );
  sg13g2_o21ai_1 _13901_ (
    .A1(addr_i_4_),
    .A2(_03766_),
    .B1(_00567_),
    .Y(_03767_)
  );
  sg13g2_nor3_1 _13902_ (
    .A(_00400_),
    .B(_00687_),
    .C(_00346_),
    .Y(_03768_)
  );
  sg13g2_a22oi_1 _13903_ (
    .A1(_00799_),
    .A2(_03767_),
    .B1(_03768_),
    .B2(_06619_),
    .Y(_03769_)
  );
  sg13g2_o21ai_1 _13904_ (
    .A1(_08564_),
    .A2(_00664_),
    .B1(_00147_),
    .Y(_03770_)
  );
  sg13g2_nand2_1 _13905_ (
    .A(_00347_),
    .B(_03770_),
    .Y(_03771_)
  );
  sg13g2_nand2_1 _13906_ (
    .A(_08520_),
    .B(_00785_),
    .Y(_03772_)
  );
  sg13g2_a21oi_1 _13907_ (
    .A1(_08852_),
    .A2(_03772_),
    .B1(addr_i_7_),
    .Y(_03773_)
  );
  sg13g2_a21o_1 _13908_ (
    .A1(_03771_),
    .A2(_03773_),
    .B1(_06684_),
    .X(_03774_)
  );
  sg13g2_nand2_1 _13909_ (
    .A(addr_i_6_),
    .B(_00725_),
    .Y(_03775_)
  );
  sg13g2_nor2_1 _13910_ (
    .A(_00034_),
    .B(_03775_),
    .Y(_03777_)
  );
  sg13g2_nand2_1 _13911_ (
    .A(_03665_),
    .B(_02141_),
    .Y(_03778_)
  );
  sg13g2_a21oi_1 _13912_ (
    .A1(_04639_),
    .A2(_03778_),
    .B1(addr_i_6_),
    .Y(_03779_)
  );
  sg13g2_o21ai_1 _13913_ (
    .A1(_03777_),
    .A2(_03779_),
    .B1(_01633_),
    .Y(_03780_)
  );
  sg13g2_o21ai_1 _13914_ (
    .A1(_03769_),
    .A2(_03774_),
    .B1(_03780_),
    .Y(_03781_)
  );
  sg13g2_o21ai_1 _13915_ (
    .A1(_03764_),
    .A2(_03781_),
    .B1(addr_i_9_),
    .Y(_03782_)
  );
  sg13g2_nand2_1 _13916_ (
    .A(addr_i_5_),
    .B(_05014_),
    .Y(_03783_)
  );
  sg13g2_a21oi_1 _13917_ (
    .A1(_01203_),
    .A2(_03783_),
    .B1(addr_i_3_),
    .Y(_03784_)
  );
  sg13g2_o21ai_1 _13918_ (
    .A1(_02622_),
    .A2(_03784_),
    .B1(_06717_),
    .Y(_03785_)
  );
  sg13g2_a21oi_1 _13919_ (
    .A1(_00250_),
    .A2(_01337_),
    .B1(_02990_),
    .Y(_03786_)
  );
  sg13g2_a22oi_1 _13920_ (
    .A1(_00168_),
    .A2(_03853_),
    .B1(_03786_),
    .B2(_00067_),
    .Y(_03788_)
  );
  sg13g2_o21ai_1 _13921_ (
    .A1(_02733_),
    .A2(_02437_),
    .B1(_01694_),
    .Y(_03789_)
  );
  sg13g2_a221oi_1 _13922_ (
    .A1(_00192_),
    .A2(_00789_),
    .B1(_03789_),
    .B2(_02063_),
    .C1(addr_i_2_),
    .Y(_03790_)
  );
  sg13g2_a21oi_1 _13923_ (
    .A1(_03785_),
    .A2(_03788_),
    .B1(_03790_),
    .Y(_03791_)
  );
  sg13g2_and2_1 _13924_ (
    .A(_01948_),
    .B(_02149_),
    .X(_03792_)
  );
  sg13g2_nor2_1 _13925_ (
    .A(addr_i_3_),
    .B(_06077_),
    .Y(_03793_)
  );
  sg13g2_nor4_1 _13926_ (
    .A(_03793_),
    .B(_00933_),
    .C(_02123_),
    .D(_03039_),
    .Y(_03794_)
  );
  sg13g2_nand4_1 _13927_ (
    .A(addr_i_4_),
    .B(_00625_),
    .C(_03792_),
    .D(_03794_),
    .Y(_03795_)
  );
  sg13g2_a21oi_1 _13928_ (
    .A1(_00749_),
    .A2(_02656_),
    .B1(_01070_),
    .Y(_03796_)
  );
  sg13g2_nor2_1 _13929_ (
    .A(_07282_),
    .B(_03796_),
    .Y(_03797_)
  );
  sg13g2_a21oi_1 _13930_ (
    .A1(_03795_),
    .A2(_03797_),
    .B1(addr_i_9_),
    .Y(_03799_)
  );
  sg13g2_o21ai_1 _13931_ (
    .A1(addr_i_8_),
    .A2(_03791_),
    .B1(_03799_),
    .Y(_03800_)
  );
  sg13g2_nand3_1 _13932_ (
    .A(addr_i_10_),
    .B(_03782_),
    .C(_03800_),
    .Y(_03801_)
  );
  sg13g2_a21o_1 _13933_ (
    .A1(_03758_),
    .A2(_03801_),
    .B1(addr_i_11_),
    .X(_03802_)
  );
  sg13g2_o21ai_1 _13934_ (
    .A1(_08487_),
    .A2(_01656_),
    .B1(_02397_),
    .Y(_03803_)
  );
  sg13g2_a21oi_1 _13935_ (
    .A1(_00582_),
    .A2(_03690_),
    .B1(_01660_),
    .Y(_03804_)
  );
  sg13g2_o21ai_1 _13936_ (
    .A1(_09494_),
    .A2(_02322_),
    .B1(_00783_),
    .Y(_03805_)
  );
  sg13g2_o21ai_1 _13937_ (
    .A1(addr_i_3_),
    .A2(_03804_),
    .B1(_03805_),
    .Y(_03806_)
  );
  sg13g2_nand2_1 _13938_ (
    .A(_01571_),
    .B(_03289_),
    .Y(_03807_)
  );
  sg13g2_a21oi_1 _13939_ (
    .A1(_02804_),
    .A2(_03807_),
    .B1(_00388_),
    .Y(_03808_)
  );
  sg13g2_a21oi_1 _13940_ (
    .A1(_02257_),
    .A2(_03806_),
    .B1(_03808_),
    .Y(_03810_)
  );
  sg13g2_nor2_1 _13941_ (
    .A(_00367_),
    .B(_06927_),
    .Y(_03811_)
  );
  sg13g2_nor3_1 _13942_ (
    .A(_00479_),
    .B(addr_i_6_),
    .C(_00297_),
    .Y(_03812_)
  );
  sg13g2_a21o_1 _13943_ (
    .A1(_05247_),
    .A2(_01653_),
    .B1(_03812_),
    .X(_03813_)
  );
  sg13g2_nand4_1 _13944_ (
    .A(addr_i_3_),
    .B(addr_i_5_),
    .C(_02012_),
    .D(_02517_),
    .Y(_03814_)
  );
  sg13g2_nand2_1 _13945_ (
    .A(_01653_),
    .B(_03250_),
    .Y(_03815_)
  );
  sg13g2_a21oi_1 _13946_ (
    .A1(_03814_),
    .A2(_03815_),
    .B1(addr_i_4_),
    .Y(_03816_)
  );
  sg13g2_a22oi_1 _13947_ (
    .A1(_01365_),
    .A2(_03813_),
    .B1(_03816_),
    .B2(addr_i_8_),
    .Y(_03817_)
  );
  sg13g2_a22oi_1 _13948_ (
    .A1(_03810_),
    .A2(_03811_),
    .B1(_03817_),
    .B2(addr_i_9_),
    .Y(_03818_)
  );
  sg13g2_a21oi_1 _13949_ (
    .A1(addr_i_9_),
    .A2(_03803_),
    .B1(_03818_),
    .Y(_03819_)
  );
  sg13g2_a21oi_1 _13950_ (
    .A1(_00248_),
    .A2(_01857_),
    .B1(_01279_),
    .Y(_03821_)
  );
  sg13g2_o21ai_1 _13951_ (
    .A1(_01508_),
    .A2(_03821_),
    .B1(_00172_),
    .Y(_03822_)
  );
  sg13g2_a21oi_1 _13952_ (
    .A1(_01343_),
    .A2(_03822_),
    .B1(_02040_),
    .Y(_03823_)
  );
  sg13g2_nor2_1 _13953_ (
    .A(_03040_),
    .B(_03823_),
    .Y(_03824_)
  );
  sg13g2_o21ai_1 _13954_ (
    .A1(addr_i_10_),
    .A2(_03819_),
    .B1(_03824_),
    .Y(_03825_)
  );
  sg13g2_nand3_1 _13955_ (
    .A(addr_i_12_),
    .B(_03802_),
    .C(_03825_),
    .Y(_03826_)
  );
  sg13g2_o21ai_1 _13956_ (
    .A1(_03627_),
    .A2(_03717_),
    .B1(_03826_),
    .Y(data_o_19_)
  );
  sg13g2_o21ai_1 _13957_ (
    .A1(_04749_),
    .A2(_00934_),
    .B1(addr_i_4_),
    .Y(_03827_)
  );
  sg13g2_nand2b_1 _13958_ (
    .A_N(_01716_),
    .B(_03827_),
    .Y(_03828_)
  );
  sg13g2_nor2_1 _13959_ (
    .A(_00543_),
    .B(_01353_),
    .Y(_03829_)
  );
  sg13g2_a22oi_1 _13960_ (
    .A1(addr_i_3_),
    .A2(_03828_),
    .B1(_03829_),
    .B2(addr_i_7_),
    .Y(_03831_)
  );
  sg13g2_o21ai_1 _13961_ (
    .A1(_02634_),
    .A2(_08852_),
    .B1(_01230_),
    .Y(_03832_)
  );
  sg13g2_nand2_1 _13962_ (
    .A(_00650_),
    .B(_09475_),
    .Y(_03833_)
  );
  sg13g2_a22oi_1 _13963_ (
    .A1(addr_i_3_),
    .A2(_03833_),
    .B1(_01746_),
    .B2(_00032_),
    .Y(_03834_)
  );
  sg13g2_a22oi_1 _13964_ (
    .A1(_00428_),
    .A2(_03832_),
    .B1(_03834_),
    .B2(addr_i_8_),
    .Y(_03835_)
  );
  sg13g2_nand2b_1 _13965_ (
    .A_N(_03831_),
    .B(_03835_),
    .Y(_03836_)
  );
  sg13g2_o21ai_1 _13966_ (
    .A1(_00269_),
    .A2(_02598_),
    .B1(_01355_),
    .Y(_03837_)
  );
  sg13g2_o21ai_1 _13967_ (
    .A1(_00746_),
    .A2(_01986_),
    .B1(_00744_),
    .Y(_03838_)
  );
  sg13g2_nand2_1 _13968_ (
    .A(_01384_),
    .B(_01084_),
    .Y(_03839_)
  );
  sg13g2_nand2_1 _13969_ (
    .A(_02462_),
    .B(_03839_),
    .Y(_03840_)
  );
  sg13g2_nand4_1 _13970_ (
    .A(addr_i_7_),
    .B(_03837_),
    .C(_03838_),
    .D(_03840_),
    .Y(_03843_)
  );
  sg13g2_a21oi_1 _13971_ (
    .A1(addr_i_6_),
    .A2(_01097_),
    .B1(addr_i_7_),
    .Y(_03844_)
  );
  sg13g2_nand2_1 _13972_ (
    .A(addr_i_2_),
    .B(_05678_),
    .Y(_03845_)
  );
  sg13g2_nor2_1 _13973_ (
    .A(_04450_),
    .B(_01539_),
    .Y(_03846_)
  );
  sg13g2_a21oi_1 _13974_ (
    .A1(_00998_),
    .A2(_03845_),
    .B1(_03846_),
    .Y(_03847_)
  );
  sg13g2_nor2_1 _13975_ (
    .A(_07492_),
    .B(_00583_),
    .Y(_03848_)
  );
  sg13g2_o21ai_1 _13976_ (
    .A1(_01222_),
    .A2(_03848_),
    .B1(addr_i_8_),
    .Y(_03849_)
  );
  sg13g2_a21oi_1 _13977_ (
    .A1(_03844_),
    .A2(_03847_),
    .B1(_03849_),
    .Y(_03850_)
  );
  sg13g2_a21oi_1 _13978_ (
    .A1(_03843_),
    .A2(_03850_),
    .B1(addr_i_9_),
    .Y(_03851_)
  );
  sg13g2_o21ai_1 _13979_ (
    .A1(_03842_),
    .A2(_00175_),
    .B1(_00479_),
    .Y(_03852_)
  );
  sg13g2_nor2_1 _13980_ (
    .A(_02503_),
    .B(_01243_),
    .Y(_03854_)
  );
  sg13g2_a21oi_1 _13981_ (
    .A1(_02343_),
    .A2(_03854_),
    .B1(_00435_),
    .Y(_03855_)
  );
  sg13g2_a21oi_1 _13982_ (
    .A1(_00442_),
    .A2(_02141_),
    .B1(_02213_),
    .Y(_03856_)
  );
  sg13g2_a221oi_1 _13983_ (
    .A1(_03852_),
    .A2(_03855_),
    .B1(_03856_),
    .B2(_02838_),
    .C1(_00112_),
    .Y(_03857_)
  );
  sg13g2_nor2_1 _13984_ (
    .A(addr_i_3_),
    .B(_02858_),
    .Y(_03858_)
  );
  sg13g2_o21ai_1 _13985_ (
    .A1(_06497_),
    .A2(_03858_),
    .B1(_00744_),
    .Y(_03859_)
  );
  sg13g2_a21oi_1 _13986_ (
    .A1(addr_i_6_),
    .A2(_00019_),
    .B1(_00342_),
    .Y(_03860_)
  );
  sg13g2_o21ai_1 _13987_ (
    .A1(_02057_),
    .A2(_03860_),
    .B1(addr_i_3_),
    .Y(_03861_)
  );
  sg13g2_nand4_1 _13988_ (
    .A(addr_i_7_),
    .B(_02187_),
    .C(_03859_),
    .D(_03861_),
    .Y(_03862_)
  );
  sg13g2_o21ai_1 _13989_ (
    .A1(addr_i_4_),
    .A2(_03637_),
    .B1(_02683_),
    .Y(_03863_)
  );
  sg13g2_nand3_1 _13990_ (
    .A(addr_i_4_),
    .B(addr_i_5_),
    .C(_00447_),
    .Y(_03865_)
  );
  sg13g2_nand3_1 _13991_ (
    .A(addr_i_3_),
    .B(_02529_),
    .C(_03865_),
    .Y(_03866_)
  );
  sg13g2_o21ai_1 _13992_ (
    .A1(addr_i_3_),
    .A2(_03863_),
    .B1(_03866_),
    .Y(_03867_)
  );
  sg13g2_o21ai_1 _13993_ (
    .A1(addr_i_2_),
    .A2(_03842_),
    .B1(addr_i_3_),
    .Y(_03868_)
  );
  sg13g2_o21ai_1 _13994_ (
    .A1(addr_i_3_),
    .A2(_03089_),
    .B1(_03868_),
    .Y(_03869_)
  );
  sg13g2_a21oi_1 _13995_ (
    .A1(_00381_),
    .A2(_03869_),
    .B1(_02294_),
    .Y(_03870_)
  );
  sg13g2_nand2_1 _13996_ (
    .A(_04086_),
    .B(_07447_),
    .Y(_03871_)
  );
  sg13g2_nand2_1 _13997_ (
    .A(_01834_),
    .B(_03871_),
    .Y(_03872_)
  );
  sg13g2_o21ai_1 _13998_ (
    .A1(addr_i_3_),
    .A2(_02928_),
    .B1(_07105_),
    .Y(_03873_)
  );
  sg13g2_o21ai_1 _13999_ (
    .A1(_03872_),
    .A2(_03873_),
    .B1(_06684_),
    .Y(_03874_)
  );
  sg13g2_a22oi_1 _14000_ (
    .A1(addr_i_7_),
    .A2(_03867_),
    .B1(_03870_),
    .B2(_03874_),
    .Y(_03876_)
  );
  sg13g2_a22oi_1 _14001_ (
    .A1(_03857_),
    .A2(_03862_),
    .B1(_03876_),
    .B2(_09315_),
    .Y(_03877_)
  );
  sg13g2_a22oi_1 _14002_ (
    .A1(_03836_),
    .A2(_03851_),
    .B1(addr_i_10_),
    .B2(_03877_),
    .Y(_03878_)
  );
  sg13g2_o21ai_1 _14003_ (
    .A1(addr_i_2_),
    .A2(_00074_),
    .B1(_07160_),
    .Y(_03879_)
  );
  sg13g2_nor2_1 _14004_ (
    .A(_00316_),
    .B(_08863_),
    .Y(_03880_)
  );
  sg13g2_a221oi_1 _14005_ (
    .A1(addr_i_4_),
    .A2(_03879_),
    .B1(_03880_),
    .B2(addr_i_2_),
    .C1(_09507_),
    .Y(_03881_)
  );
  sg13g2_nand3_1 _14006_ (
    .A(addr_i_4_),
    .B(addr_i_5_),
    .C(_02558_),
    .Y(_03882_)
  );
  sg13g2_o21ai_1 _14007_ (
    .A1(_04494_),
    .A2(_01570_),
    .B1(_03882_),
    .Y(_03883_)
  );
  sg13g2_a221oi_1 _14008_ (
    .A1(_01215_),
    .A2(_01338_),
    .B1(_03883_),
    .B2(addr_i_2_),
    .C1(_02105_),
    .Y(_03884_)
  );
  sg13g2_a21o_1 _14009_ (
    .A1(_02271_),
    .A2(_03881_),
    .B1(_03884_),
    .X(_03885_)
  );
  sg13g2_a21oi_1 _14010_ (
    .A1(_01384_),
    .A2(_01084_),
    .B1(addr_i_3_),
    .Y(_03887_)
  );
  sg13g2_o21ai_1 _14011_ (
    .A1(_01375_),
    .A2(_03887_),
    .B1(addr_i_6_),
    .Y(_03888_)
  );
  sg13g2_nand3_1 _14012_ (
    .A(_03374_),
    .B(_02187_),
    .C(_03888_),
    .Y(_03889_)
  );
  sg13g2_nor2_1 _14013_ (
    .A(addr_i_7_),
    .B(_01610_),
    .Y(_03890_)
  );
  sg13g2_nand3_1 _14014_ (
    .A(_01652_),
    .B(_03167_),
    .C(_01029_),
    .Y(_03891_)
  );
  sg13g2_nor2_1 _14015_ (
    .A(_02086_),
    .B(_01264_),
    .Y(_03892_)
  );
  sg13g2_o21ai_1 _14016_ (
    .A1(_02441_),
    .A2(_03892_),
    .B1(addr_i_5_),
    .Y(_03893_)
  );
  sg13g2_nand4_1 _14017_ (
    .A(_02930_),
    .B(_03890_),
    .C(_03891_),
    .D(_03893_),
    .Y(_03894_)
  );
  sg13g2_nand3_1 _14018_ (
    .A(addr_i_10_),
    .B(_03889_),
    .C(_03894_),
    .Y(_03895_)
  );
  sg13g2_a21oi_1 _14019_ (
    .A1(_00423_),
    .A2(_03885_),
    .B1(_03895_),
    .Y(_03896_)
  );
  sg13g2_or2_1 _14020_ (
    .A(_03878_),
    .B(_03896_),
    .X(_03898_)
  );
  sg13g2_nor2_1 _14021_ (
    .A(addr_i_3_),
    .B(_01635_),
    .Y(_03899_)
  );
  sg13g2_nor2_1 _14022_ (
    .A(_02264_),
    .B(_03899_),
    .Y(_03900_)
  );
  sg13g2_a22oi_1 _14023_ (
    .A1(_00347_),
    .A2(_02184_),
    .B1(_00369_),
    .B2(addr_i_2_),
    .Y(_03901_)
  );
  sg13g2_a21oi_1 _14024_ (
    .A1(addr_i_2_),
    .A2(_03900_),
    .B1(_03901_),
    .Y(_03902_)
  );
  sg13g2_nor2_1 _14025_ (
    .A(addr_i_3_),
    .B(_08763_),
    .Y(_03903_)
  );
  sg13g2_o21ai_1 _14026_ (
    .A1(_03501_),
    .A2(_03903_),
    .B1(_00293_),
    .Y(_03904_)
  );
  sg13g2_a21oi_1 _14027_ (
    .A1(addr_i_2_),
    .A2(addr_i_6_),
    .B1(addr_i_5_),
    .Y(_03905_)
  );
  sg13g2_nor2_1 _14028_ (
    .A(_00342_),
    .B(_03905_),
    .Y(_03906_)
  );
  sg13g2_o21ai_1 _14029_ (
    .A1(_09348_),
    .A2(_03906_),
    .B1(addr_i_3_),
    .Y(_03907_)
  );
  sg13g2_nand4_1 _14030_ (
    .A(_00429_),
    .B(_00907_),
    .C(_03904_),
    .D(_03907_),
    .Y(_03909_)
  );
  sg13g2_o21ai_1 _14031_ (
    .A1(_01099_),
    .A2(_03902_),
    .B1(_03909_),
    .Y(_03910_)
  );
  sg13g2_o21ai_1 _14032_ (
    .A1(_05236_),
    .A2(_00095_),
    .B1(addr_i_5_),
    .Y(_03911_)
  );
  sg13g2_a21oi_1 _14033_ (
    .A1(_02623_),
    .A2(_07967_),
    .B1(addr_i_3_),
    .Y(_03912_)
  );
  sg13g2_nand2_1 _14034_ (
    .A(_03911_),
    .B(_03912_),
    .Y(_03913_)
  );
  sg13g2_nor2_1 _14035_ (
    .A(addr_i_4_),
    .B(_01592_),
    .Y(_03914_)
  );
  sg13g2_nor2_1 _14036_ (
    .A(_04550_),
    .B(_08089_),
    .Y(_03915_)
  );
  sg13g2_nor2_1 _14037_ (
    .A(_00637_),
    .B(_03915_),
    .Y(_03916_)
  );
  sg13g2_nor4_1 _14038_ (
    .A(_06364_),
    .B(_00624_),
    .C(_03914_),
    .D(_03916_),
    .Y(_03917_)
  );
  sg13g2_a21oi_1 _14039_ (
    .A1(_00019_),
    .A2(_00994_),
    .B1(addr_i_4_),
    .Y(_03918_)
  );
  sg13g2_nor3_1 _14040_ (
    .A(addr_i_6_),
    .B(_00632_),
    .C(_03918_),
    .Y(_03920_)
  );
  sg13g2_o21ai_1 _14041_ (
    .A1(_03917_),
    .A2(_03920_),
    .B1(addr_i_3_),
    .Y(_03921_)
  );
  sg13g2_nor2_1 _14042_ (
    .A(_07967_),
    .B(_03566_),
    .Y(_03922_)
  );
  sg13g2_o21ai_1 _14043_ (
    .A1(_00961_),
    .A2(_03922_),
    .B1(_02683_),
    .Y(_03923_)
  );
  sg13g2_a221oi_1 _14044_ (
    .A1(_03913_),
    .A2(_03921_),
    .B1(_03923_),
    .B2(_03263_),
    .C1(_03617_),
    .Y(_03924_)
  );
  sg13g2_o21ai_1 _14045_ (
    .A1(_03910_),
    .A2(_03924_),
    .B1(_05203_),
    .Y(_03925_)
  );
  sg13g2_and2_1 _14046_ (
    .A(addr_i_11_),
    .B(_03925_),
    .X(_03926_)
  );
  sg13g2_nand2_1 _14047_ (
    .A(_08166_),
    .B(_01014_),
    .Y(_03927_)
  );
  sg13g2_nand2_1 _14048_ (
    .A(_00339_),
    .B(_03927_),
    .Y(_03928_)
  );
  sg13g2_a21oi_1 _14049_ (
    .A1(_01265_),
    .A2(_01715_),
    .B1(_04461_),
    .Y(_03929_)
  );
  sg13g2_a22oi_1 _14050_ (
    .A1(_00910_),
    .A2(_03928_),
    .B1(_03929_),
    .B2(_02055_),
    .Y(_03931_)
  );
  sg13g2_nand2_1 _14051_ (
    .A(_02020_),
    .B(_01406_),
    .Y(_03932_)
  );
  sg13g2_a22oi_1 _14052_ (
    .A1(addr_i_3_),
    .A2(_03932_),
    .B1(_00206_),
    .B2(_00351_),
    .Y(_03933_)
  );
  sg13g2_a21oi_1 _14053_ (
    .A1(_01475_),
    .A2(_03931_),
    .B1(_03933_),
    .Y(_03934_)
  );
  sg13g2_o21ai_1 _14054_ (
    .A1(_07558_),
    .A2(_07724_),
    .B1(addr_i_8_),
    .Y(_03935_)
  );
  sg13g2_nand2_1 _14055_ (
    .A(addr_i_2_),
    .B(_03167_),
    .Y(_03936_)
  );
  sg13g2_nand2_1 _14056_ (
    .A(_04650_),
    .B(_00371_),
    .Y(_03937_)
  );
  sg13g2_a21oi_1 _14057_ (
    .A1(_01160_),
    .A2(_02898_),
    .B1(addr_i_3_),
    .Y(_03938_)
  );
  sg13g2_a22oi_1 _14058_ (
    .A1(_00607_),
    .A2(_03936_),
    .B1(_03937_),
    .B2(_03938_),
    .Y(_03939_)
  );
  sg13g2_nand2_1 _14059_ (
    .A(_00531_),
    .B(_00719_),
    .Y(_03940_)
  );
  sg13g2_o21ai_1 _14060_ (
    .A1(addr_i_2_),
    .A2(addr_i_6_),
    .B1(addr_i_4_),
    .Y(_03942_)
  );
  sg13g2_nand2_1 _14061_ (
    .A(addr_i_3_),
    .B(_03942_),
    .Y(_03943_)
  );
  sg13g2_nand2b_1 _14062_ (
    .A_N(_03942_),
    .B(_00347_),
    .Y(_03944_)
  );
  sg13g2_a21oi_1 _14063_ (
    .A1(_03943_),
    .A2(_03944_),
    .B1(addr_i_5_),
    .Y(_03945_)
  );
  sg13g2_a22oi_1 _14064_ (
    .A1(_01216_),
    .A2(_03940_),
    .B1(_03945_),
    .B2(_00600_),
    .Y(_03946_)
  );
  sg13g2_a21oi_1 _14065_ (
    .A1(_02263_),
    .A2(_03939_),
    .B1(_03946_),
    .Y(_03947_)
  );
  sg13g2_o21ai_1 _14066_ (
    .A1(_03934_),
    .A2(_03935_),
    .B1(_03947_),
    .Y(_03948_)
  );
  sg13g2_a22oi_1 _14067_ (
    .A1(addr_i_3_),
    .A2(_02585_),
    .B1(_00746_),
    .B2(_02598_),
    .Y(_03949_)
  );
  sg13g2_a22oi_1 _14068_ (
    .A1(_00065_),
    .A2(_02329_),
    .B1(_01091_),
    .B2(addr_i_7_),
    .Y(_03950_)
  );
  sg13g2_o21ai_1 _14069_ (
    .A1(addr_i_4_),
    .A2(_03949_),
    .B1(_03950_),
    .Y(_03951_)
  );
  sg13g2_nand2_1 _14070_ (
    .A(addr_i_5_),
    .B(_00711_),
    .Y(_03954_)
  );
  sg13g2_nand3_1 _14071_ (
    .A(_00428_),
    .B(_09476_),
    .C(_03954_),
    .Y(_03955_)
  );
  sg13g2_nand3_1 _14072_ (
    .A(_09061_),
    .B(_02854_),
    .C(_03428_),
    .Y(_03956_)
  );
  sg13g2_nand4_1 _14073_ (
    .A(addr_i_8_),
    .B(_03951_),
    .C(_03955_),
    .D(_03956_),
    .Y(_03957_)
  );
  sg13g2_o21ai_1 _14074_ (
    .A1(_05722_),
    .A2(_07746_),
    .B1(addr_i_3_),
    .Y(_03958_)
  );
  sg13g2_nand2b_1 _14075_ (
    .A_N(_01192_),
    .B(_03958_),
    .Y(_03959_)
  );
  sg13g2_o21ai_1 _14076_ (
    .A1(_00586_),
    .A2(_03842_),
    .B1(_00380_),
    .Y(_03960_)
  );
  sg13g2_a221oi_1 _14077_ (
    .A1(addr_i_2_),
    .A2(_03959_),
    .B1(_03960_),
    .B2(_03809_),
    .C1(addr_i_6_),
    .Y(_03961_)
  );
  sg13g2_nor2_1 _14078_ (
    .A(_04362_),
    .B(_04218_),
    .Y(_03962_)
  );
  sg13g2_nor2_1 _14079_ (
    .A(addr_i_4_),
    .B(_02843_),
    .Y(_03963_)
  );
  sg13g2_a22oi_1 _14080_ (
    .A1(_02496_),
    .A2(_03962_),
    .B1(_03963_),
    .B2(_00006_),
    .Y(_03965_)
  );
  sg13g2_nor3_1 _14081_ (
    .A(_09497_),
    .B(_00021_),
    .C(_03033_),
    .Y(_03966_)
  );
  sg13g2_or4_1 _14082_ (
    .A(addr_i_8_),
    .B(_03961_),
    .C(_03965_),
    .D(_03966_),
    .X(_03967_)
  );
  sg13g2_nand2_1 _14083_ (
    .A(_03957_),
    .B(_03967_),
    .Y(_03968_)
  );
  sg13g2_nand2_1 _14084_ (
    .A(_00319_),
    .B(_00591_),
    .Y(_03969_)
  );
  sg13g2_nor2_1 _14085_ (
    .A(_09038_),
    .B(_00577_),
    .Y(_03970_)
  );
  sg13g2_o21ai_1 _14086_ (
    .A1(_00346_),
    .A2(_03970_),
    .B1(addr_i_2_),
    .Y(_03971_)
  );
  sg13g2_a21o_1 _14087_ (
    .A1(_03969_),
    .A2(_03971_),
    .B1(_02064_),
    .X(_03972_)
  );
  sg13g2_a21oi_1 _14088_ (
    .A1(_00435_),
    .A2(_00079_),
    .B1(_00483_),
    .Y(_03973_)
  );
  sg13g2_o21ai_1 _14089_ (
    .A1(_08089_),
    .A2(_01022_),
    .B1(_05281_),
    .Y(_03974_)
  );
  sg13g2_nand3_1 _14090_ (
    .A(_01658_),
    .B(_02156_),
    .C(_03974_),
    .Y(_03976_)
  );
  sg13g2_o21ai_1 _14091_ (
    .A1(_03973_),
    .A2(_03976_),
    .B1(addr_i_5_),
    .Y(_03977_)
  );
  sg13g2_nand3_1 _14092_ (
    .A(_03746_),
    .B(_03972_),
    .C(_03977_),
    .Y(_03978_)
  );
  sg13g2_nand2_1 _14093_ (
    .A(_00357_),
    .B(_02001_),
    .Y(_03979_)
  );
  sg13g2_nor2_1 _14094_ (
    .A(addr_i_4_),
    .B(_01066_),
    .Y(_03980_)
  );
  sg13g2_a21o_1 _14095_ (
    .A1(addr_i_4_),
    .A2(_03979_),
    .B1(_03980_),
    .X(_03981_)
  );
  sg13g2_a221oi_1 _14096_ (
    .A1(_01450_),
    .A2(_02948_),
    .B1(_03981_),
    .B2(_00949_),
    .C1(_01285_),
    .Y(_03982_)
  );
  sg13g2_o21ai_1 _14097_ (
    .A1(_03759_),
    .A2(_00824_),
    .B1(_00648_),
    .Y(_03983_)
  );
  sg13g2_a22oi_1 _14098_ (
    .A1(addr_i_2_),
    .A2(_04418_),
    .B1(_03676_),
    .B2(addr_i_3_),
    .Y(_03984_)
  );
  sg13g2_nor3_1 _14099_ (
    .A(_00593_),
    .B(_03270_),
    .C(_03172_),
    .Y(_03985_)
  );
  sg13g2_o21ai_1 _14100_ (
    .A1(_03984_),
    .A2(_03985_),
    .B1(addr_i_4_),
    .Y(_03987_)
  );
  sg13g2_nand4_1 _14101_ (
    .A(_01310_),
    .B(_00131_),
    .C(_03983_),
    .D(_03987_),
    .Y(_03988_)
  );
  sg13g2_nand2_1 _14102_ (
    .A(_00385_),
    .B(_03988_),
    .Y(_03989_)
  );
  sg13g2_a22oi_1 _14103_ (
    .A1(_01043_),
    .A2(_03978_),
    .B1(_03982_),
    .B2(_03989_),
    .Y(_03990_)
  );
  sg13g2_a22oi_1 _14104_ (
    .A1(addr_i_9_),
    .A2(_03968_),
    .B1(_03990_),
    .B2(addr_i_10_),
    .Y(_03991_)
  );
  sg13g2_a22oi_1 _14105_ (
    .A1(_01174_),
    .A2(_03948_),
    .B1(_03991_),
    .B2(addr_i_11_),
    .Y(_03992_)
  );
  sg13g2_buf_1 _14106_ (
    .A(_05943_),
    .X(_03993_)
  );
  sg13g2_o21ai_1 _14107_ (
    .A1(_03993_),
    .A2(_06740_),
    .B1(_00561_),
    .Y(_03994_)
  );
  sg13g2_o21ai_1 _14108_ (
    .A1(_00184_),
    .A2(_00789_),
    .B1(_03994_),
    .Y(_03995_)
  );
  sg13g2_nand3_1 _14109_ (
    .A(addr_i_2_),
    .B(_06895_),
    .C(_01007_),
    .Y(_03996_)
  );
  sg13g2_nor2_1 _14110_ (
    .A(_01517_),
    .B(_08807_),
    .Y(_03998_)
  );
  sg13g2_o21ai_1 _14111_ (
    .A1(addr_i_3_),
    .A2(_00990_),
    .B1(_01007_),
    .Y(_03999_)
  );
  sg13g2_a22oi_1 _14112_ (
    .A1(addr_i_2_),
    .A2(_03999_),
    .B1(_02269_),
    .B2(addr_i_7_),
    .Y(_04000_)
  );
  sg13g2_a22oi_1 _14113_ (
    .A1(_03996_),
    .A2(_03998_),
    .B1(_04000_),
    .B2(_00084_),
    .Y(_04001_)
  );
  sg13g2_a22oi_1 _14114_ (
    .A1(_01630_),
    .A2(_03995_),
    .B1(_04001_),
    .B2(_03259_),
    .Y(_04002_)
  );
  sg13g2_a21oi_1 _14115_ (
    .A1(_00069_),
    .A2(_00055_),
    .B1(_02105_),
    .Y(_04003_)
  );
  sg13g2_o21ai_1 _14116_ (
    .A1(_02848_),
    .A2(_04003_),
    .B1(addr_i_2_),
    .Y(_04004_)
  );
  sg13g2_nand2b_1 _14117_ (
    .A_N(_03589_),
    .B(_04004_),
    .Y(_04005_)
  );
  sg13g2_nor2_1 _14118_ (
    .A(_00334_),
    .B(_03153_),
    .Y(_04006_)
  );
  sg13g2_a22oi_1 _14119_ (
    .A1(_00492_),
    .A2(_02742_),
    .B1(_02154_),
    .B2(addr_i_2_),
    .Y(_04007_)
  );
  sg13g2_a22oi_1 _14120_ (
    .A1(addr_i_2_),
    .A2(_04006_),
    .B1(_04007_),
    .B2(_00084_),
    .Y(_04009_)
  );
  sg13g2_o21ai_1 _14121_ (
    .A1(_02191_),
    .A2(_01193_),
    .B1(_00782_),
    .Y(_04010_)
  );
  sg13g2_a22oi_1 _14122_ (
    .A1(_00172_),
    .A2(_04005_),
    .B1(_04009_),
    .B2(_04010_),
    .Y(_04011_)
  );
  sg13g2_o21ai_1 _14123_ (
    .A1(_04002_),
    .A2(_04011_),
    .B1(_05214_),
    .Y(_04012_)
  );
  sg13g2_a221oi_1 _14124_ (
    .A1(_03898_),
    .A2(_03926_),
    .B1(_03992_),
    .B2(_04012_),
    .C1(addr_i_12_),
    .Y(_04013_)
  );
  sg13g2_a21oi_1 _14125_ (
    .A1(addr_i_7_),
    .A2(_00150_),
    .B1(addr_i_4_),
    .Y(_04014_)
  );
  sg13g2_a22oi_1 _14126_ (
    .A1(addr_i_4_),
    .A2(_01128_),
    .B1(_04014_),
    .B2(addr_i_3_),
    .Y(_04015_)
  );
  sg13g2_nor2_1 _14127_ (
    .A(_00001_),
    .B(_00632_),
    .Y(_04016_)
  );
  sg13g2_a22oi_1 _14128_ (
    .A1(addr_i_4_),
    .A2(_04016_),
    .B1(_00683_),
    .B2(_01935_),
    .Y(_04017_)
  );
  sg13g2_a22oi_1 _14129_ (
    .A1(_05833_),
    .A2(_01216_),
    .B1(_04015_),
    .B2(_04017_),
    .Y(_04018_)
  );
  sg13g2_nor2_1 _14130_ (
    .A(_00617_),
    .B(_01202_),
    .Y(_04020_)
  );
  sg13g2_o21ai_1 _14131_ (
    .A1(addr_i_3_),
    .A2(_02850_),
    .B1(_04020_),
    .Y(_04021_)
  );
  sg13g2_nand2_1 _14132_ (
    .A(_00024_),
    .B(_00650_),
    .Y(_04022_)
  );
  sg13g2_a22oi_1 _14133_ (
    .A1(addr_i_3_),
    .A2(_04022_),
    .B1(_00133_),
    .B2(_00053_),
    .Y(_04023_)
  );
  sg13g2_a22oi_1 _14134_ (
    .A1(_09487_),
    .A2(_04021_),
    .B1(_04023_),
    .B2(addr_i_8_),
    .Y(_04024_)
  );
  sg13g2_o21ai_1 _14135_ (
    .A1(addr_i_6_),
    .A2(_04018_),
    .B1(_04024_),
    .Y(_04025_)
  );
  sg13g2_a21oi_1 _14136_ (
    .A1(_00400_),
    .A2(_02395_),
    .B1(_02333_),
    .Y(_04026_)
  );
  sg13g2_o21ai_1 _14137_ (
    .A1(_02086_),
    .A2(_00664_),
    .B1(_01037_),
    .Y(_04027_)
  );
  sg13g2_a22oi_1 _14138_ (
    .A1(addr_i_2_),
    .A2(_04027_),
    .B1(_02143_),
    .B2(addr_i_7_),
    .Y(_04028_)
  );
  sg13g2_o21ai_1 _14139_ (
    .A1(addr_i_2_),
    .A2(_04026_),
    .B1(_04028_),
    .Y(_04029_)
  );
  sg13g2_nor2_1 _14140_ (
    .A(_00052_),
    .B(_00850_),
    .Y(_04031_)
  );
  sg13g2_o21ai_1 _14141_ (
    .A1(addr_i_3_),
    .A2(_02560_),
    .B1(_04031_),
    .Y(_04032_)
  );
  sg13g2_o21ai_1 _14142_ (
    .A1(_01881_),
    .A2(_02304_),
    .B1(_00262_),
    .Y(_04033_)
  );
  sg13g2_nand4_1 _14143_ (
    .A(addr_i_8_),
    .B(_04029_),
    .C(_04032_),
    .D(_04033_),
    .Y(_04034_)
  );
  sg13g2_and2_1 _14144_ (
    .A(_05203_),
    .B(_04034_),
    .X(_04035_)
  );
  sg13g2_nand2_1 _14145_ (
    .A(addr_i_10_),
    .B(_02604_),
    .Y(_04036_)
  );
  sg13g2_nor2_1 _14146_ (
    .A(_09509_),
    .B(_01954_),
    .Y(_04037_)
  );
  sg13g2_a21oi_1 _14147_ (
    .A1(addr_i_3_),
    .A2(_01645_),
    .B1(_04037_),
    .Y(_04038_)
  );
  sg13g2_nor2_1 _14148_ (
    .A(_06717_),
    .B(_04038_),
    .Y(_04039_)
  );
  sg13g2_a21oi_1 _14149_ (
    .A1(_01262_),
    .A2(_00157_),
    .B1(_04039_),
    .Y(_04040_)
  );
  sg13g2_o21ai_1 _14150_ (
    .A1(_00354_),
    .A2(_03110_),
    .B1(_00863_),
    .Y(_04042_)
  );
  sg13g2_o21ai_1 _14151_ (
    .A1(_01867_),
    .A2(_00132_),
    .B1(addr_i_5_),
    .Y(_04043_)
  );
  sg13g2_nand2b_1 _14152_ (
    .A_N(_03692_),
    .B(_04043_),
    .Y(_04044_)
  );
  sg13g2_a221oi_1 _14153_ (
    .A1(_01747_),
    .A2(_04042_),
    .B1(_04044_),
    .B2(addr_i_3_),
    .C1(addr_i_2_),
    .Y(_04045_)
  );
  sg13g2_a21oi_1 _14154_ (
    .A1(addr_i_2_),
    .A2(_04040_),
    .B1(_04045_),
    .Y(_04046_)
  );
  sg13g2_a22oi_1 _14155_ (
    .A1(_00073_),
    .A2(_00898_),
    .B1(_04036_),
    .B2(_04046_),
    .Y(_04047_)
  );
  sg13g2_nor2_1 _14156_ (
    .A(addr_i_6_),
    .B(_00454_),
    .Y(_04048_)
  );
  sg13g2_a21oi_1 _14157_ (
    .A1(_01585_),
    .A2(_01954_),
    .B1(_08188_),
    .Y(_04049_)
  );
  sg13g2_o21ai_1 _14158_ (
    .A1(addr_i_3_),
    .A2(_04048_),
    .B1(_04049_),
    .Y(_04050_)
  );
  sg13g2_a21oi_1 _14159_ (
    .A1(_00492_),
    .A2(_00434_),
    .B1(_01144_),
    .Y(_04051_)
  );
  sg13g2_a22oi_1 _14160_ (
    .A1(_08011_),
    .A2(_04050_),
    .B1(_04051_),
    .B2(addr_i_4_),
    .Y(_04053_)
  );
  sg13g2_a21o_1 _14161_ (
    .A1(addr_i_3_),
    .A2(_02090_),
    .B1(_09507_),
    .X(_04054_)
  );
  sg13g2_a21oi_1 _14162_ (
    .A1(_07558_),
    .A2(_00951_),
    .B1(_06895_),
    .Y(_04055_)
  );
  sg13g2_a22oi_1 _14163_ (
    .A1(addr_i_2_),
    .A2(_04054_),
    .B1(_04055_),
    .B2(_01794_),
    .Y(_04056_)
  );
  sg13g2_o21ai_1 _14164_ (
    .A1(_04053_),
    .A2(_04056_),
    .B1(_00215_),
    .Y(_04057_)
  );
  sg13g2_nand2_1 _14165_ (
    .A(_03029_),
    .B(_04057_),
    .Y(_04058_)
  );
  sg13g2_a22oi_1 _14166_ (
    .A1(_04025_),
    .A2(_04035_),
    .B1(_04047_),
    .B2(_04058_),
    .Y(_04059_)
  );
  sg13g2_nor2_1 _14167_ (
    .A(_08741_),
    .B(_04837_),
    .Y(_04060_)
  );
  sg13g2_and2_1 _14168_ (
    .A(_02489_),
    .B(_04060_),
    .X(_04061_)
  );
  sg13g2_nor2_1 _14169_ (
    .A(_02777_),
    .B(_01305_),
    .Y(_04062_)
  );
  sg13g2_a22oi_1 _14170_ (
    .A1(_01095_),
    .A2(_02057_),
    .B1(_04062_),
    .B2(addr_i_3_),
    .Y(_04065_)
  );
  sg13g2_o21ai_1 _14171_ (
    .A1(_04061_),
    .A2(_04065_),
    .B1(_01861_),
    .Y(_04066_)
  );
  sg13g2_nand2_1 _14172_ (
    .A(_00020_),
    .B(_00442_),
    .Y(_04067_)
  );
  sg13g2_buf_1 _14173_ (
    .A(_03809_),
    .X(_04068_)
  );
  sg13g2_a21oi_1 _14174_ (
    .A1(_04067_),
    .A2(_03189_),
    .B1(_04068_),
    .Y(_04069_)
  );
  sg13g2_nor2_1 _14175_ (
    .A(_07248_),
    .B(_02327_),
    .Y(_04070_)
  );
  sg13g2_nor2_1 _14176_ (
    .A(_00697_),
    .B(_04070_),
    .Y(_04071_)
  );
  sg13g2_o21ai_1 _14177_ (
    .A1(_04069_),
    .A2(_04071_),
    .B1(addr_i_6_),
    .Y(_04072_)
  );
  sg13g2_nand3_1 _14178_ (
    .A(_03953_),
    .B(_00021_),
    .C(_08111_),
    .Y(_04073_)
  );
  sg13g2_a21oi_1 _14179_ (
    .A1(_02987_),
    .A2(_04073_),
    .B1(_02344_),
    .Y(_04074_)
  );
  sg13g2_a22oi_1 _14180_ (
    .A1(_00223_),
    .A2(_03572_),
    .B1(_04074_),
    .B2(addr_i_8_),
    .Y(_04076_)
  );
  sg13g2_a21o_1 _14181_ (
    .A1(addr_i_6_),
    .A2(addr_i_5_),
    .B1(addr_i_4_),
    .X(_04077_)
  );
  sg13g2_a21oi_1 _14182_ (
    .A1(_08431_),
    .A2(_04077_),
    .B1(_00697_),
    .Y(_04078_)
  );
  sg13g2_a22oi_1 _14183_ (
    .A1(_01020_),
    .A2(_01309_),
    .B1(_04078_),
    .B2(_00290_),
    .Y(_04079_)
  );
  sg13g2_a22oi_1 _14184_ (
    .A1(_04072_),
    .A2(_04076_),
    .B1(addr_i_9_),
    .B2(_04079_),
    .Y(_04080_)
  );
  sg13g2_a21oi_1 _14185_ (
    .A1(_04066_),
    .A2(_04080_),
    .B1(addr_i_10_),
    .Y(_04081_)
  );
  sg13g2_a21oi_1 _14186_ (
    .A1(_00441_),
    .A2(_03540_),
    .B1(addr_i_4_),
    .Y(_04082_)
  );
  sg13g2_o21ai_1 _14187_ (
    .A1(_04483_),
    .A2(_04082_),
    .B1(addr_i_6_),
    .Y(_04083_)
  );
  sg13g2_o21ai_1 _14188_ (
    .A1(addr_i_7_),
    .A2(_05258_),
    .B1(addr_i_4_),
    .Y(_04084_)
  );
  sg13g2_nand2b_1 _14189_ (
    .A_N(_03918_),
    .B(_04084_),
    .Y(_04085_)
  );
  sg13g2_nand2_1 _14190_ (
    .A(addr_i_4_),
    .B(_06729_),
    .Y(_04087_)
  );
  sg13g2_a21oi_1 _14191_ (
    .A1(_04087_),
    .A2(_01343_),
    .B1(addr_i_5_),
    .Y(_04088_)
  );
  sg13g2_a22oi_1 _14192_ (
    .A1(_00388_),
    .A2(_04085_),
    .B1(_04088_),
    .B2(_00116_),
    .Y(_04089_)
  );
  sg13g2_a21oi_1 _14193_ (
    .A1(_02942_),
    .A2(_04083_),
    .B1(_04089_),
    .Y(_04090_)
  );
  sg13g2_nand2_1 _14194_ (
    .A(addr_i_4_),
    .B(_00140_),
    .Y(_04091_)
  );
  sg13g2_nand2_1 _14195_ (
    .A(addr_i_6_),
    .B(_00462_),
    .Y(_04092_)
  );
  sg13g2_nand2_1 _14196_ (
    .A(_00593_),
    .B(_04092_),
    .Y(_04093_)
  );
  sg13g2_nand3_1 _14197_ (
    .A(_01715_),
    .B(_04091_),
    .C(_04093_),
    .Y(_04094_)
  );
  sg13g2_nand2_1 _14198_ (
    .A(addr_i_3_),
    .B(_03842_),
    .Y(_04095_)
  );
  sg13g2_nand2_1 _14199_ (
    .A(_02501_),
    .B(_04095_),
    .Y(_04096_)
  );
  sg13g2_a21oi_1 _14200_ (
    .A1(_00104_),
    .A2(_00228_),
    .B1(addr_i_3_),
    .Y(_04098_)
  );
  sg13g2_nor3_1 _14201_ (
    .A(_04981_),
    .B(_00840_),
    .C(_00244_),
    .Y(_04099_)
  );
  sg13g2_o21ai_1 _14202_ (
    .A1(_03853_),
    .A2(_04099_),
    .B1(_02498_),
    .Y(_04100_)
  );
  sg13g2_o21ai_1 _14203_ (
    .A1(_04096_),
    .A2(_04098_),
    .B1(_04100_),
    .Y(_04101_)
  );
  sg13g2_a22oi_1 _14204_ (
    .A1(_01119_),
    .A2(_04094_),
    .B1(_04101_),
    .B2(_01351_),
    .Y(_04102_)
  );
  sg13g2_o21ai_1 _14205_ (
    .A1(addr_i_8_),
    .A2(_04090_),
    .B1(_04102_),
    .Y(_04103_)
  );
  sg13g2_nand2_1 _14206_ (
    .A(_04081_),
    .B(_04103_),
    .Y(_04104_)
  );
  sg13g2_a21oi_1 _14207_ (
    .A1(_01892_),
    .A2(_01365_),
    .B1(_02542_),
    .Y(_04105_)
  );
  sg13g2_o21ai_1 _14208_ (
    .A1(addr_i_3_),
    .A2(_04105_),
    .B1(_02136_),
    .Y(_04106_)
  );
  sg13g2_o21ai_1 _14209_ (
    .A1(addr_i_4_),
    .A2(_08487_),
    .B1(_01668_),
    .Y(_04107_)
  );
  sg13g2_o21ai_1 _14210_ (
    .A1(_06950_),
    .A2(_03523_),
    .B1(addr_i_2_),
    .Y(_04109_)
  );
  sg13g2_nand2_1 _14211_ (
    .A(_02411_),
    .B(_04109_),
    .Y(_04110_)
  );
  sg13g2_o21ai_1 _14212_ (
    .A1(_01436_),
    .A2(_03501_),
    .B1(addr_i_5_),
    .Y(_04111_)
  );
  sg13g2_a21oi_1 _14213_ (
    .A1(_01224_),
    .A2(_04111_),
    .B1(addr_i_7_),
    .Y(_04112_)
  );
  sg13g2_o21ai_1 _14214_ (
    .A1(_04110_),
    .A2(_04112_),
    .B1(addr_i_3_),
    .Y(_04113_)
  );
  sg13g2_nand2_1 _14215_ (
    .A(addr_i_6_),
    .B(_08564_),
    .Y(_04114_)
  );
  sg13g2_a22oi_1 _14216_ (
    .A1(addr_i_7_),
    .A2(_04114_),
    .B1(_09499_),
    .B2(addr_i_3_),
    .Y(_04115_)
  );
  sg13g2_a21oi_1 _14217_ (
    .A1(_04111_),
    .A2(_04115_),
    .B1(addr_i_8_),
    .Y(_04116_)
  );
  sg13g2_o21ai_1 _14218_ (
    .A1(addr_i_7_),
    .A2(_03033_),
    .B1(_01277_),
    .Y(_04117_)
  );
  sg13g2_nand3_1 _14219_ (
    .A(addr_i_8_),
    .B(_01199_),
    .C(_04117_),
    .Y(_04118_)
  );
  sg13g2_o21ai_1 _14220_ (
    .A1(addr_i_5_),
    .A2(_02462_),
    .B1(addr_i_2_),
    .Y(_04120_)
  );
  sg13g2_and2_1 _14221_ (
    .A(addr_i_3_),
    .B(_00591_),
    .X(_04121_)
  );
  sg13g2_nor2b_1 _14222_ (
    .A(_04121_),
    .B_N(_02850_),
    .Y(_04122_)
  );
  sg13g2_a22oi_1 _14223_ (
    .A1(addr_i_4_),
    .A2(_04120_),
    .B1(_04122_),
    .B2(addr_i_7_),
    .Y(_04123_)
  );
  sg13g2_nor2_1 _14224_ (
    .A(_04118_),
    .B(_04123_),
    .Y(_04124_)
  );
  sg13g2_a22oi_1 _14225_ (
    .A1(_04113_),
    .A2(_04116_),
    .B1(addr_i_9_),
    .B2(_04124_),
    .Y(_04125_)
  );
  sg13g2_a22oi_1 _14226_ (
    .A1(addr_i_9_),
    .A2(_04107_),
    .B1(_04125_),
    .B2(addr_i_10_),
    .Y(_04126_)
  );
  sg13g2_a22oi_1 _14227_ (
    .A1(_01350_),
    .A2(_04106_),
    .B1(_04126_),
    .B2(_01640_),
    .Y(_04127_)
  );
  sg13g2_a22oi_1 _14228_ (
    .A1(_04059_),
    .A2(_04104_),
    .B1(_00812_),
    .B2(_04127_),
    .Y(_04128_)
  );
  sg13g2_or2_1 _14229_ (
    .A(_04013_),
    .B(_04128_),
    .X(data_o_1_)
  );
  sg13g2_nor2_1 _14230_ (
    .A(_02525_),
    .B(_02207_),
    .Y(_04130_)
  );
  sg13g2_nor2_1 _14231_ (
    .A(addr_i_7_),
    .B(_01355_),
    .Y(_04131_)
  );
  sg13g2_a21oi_1 _14232_ (
    .A1(_01892_),
    .A2(_04130_),
    .B1(_04131_),
    .Y(_04132_)
  );
  sg13g2_o21ai_1 _14233_ (
    .A1(_02040_),
    .A2(_04132_),
    .B1(addr_i_11_),
    .Y(_04133_)
  );
  sg13g2_a21oi_1 _14234_ (
    .A1(_00831_),
    .A2(_00173_),
    .B1(addr_i_3_),
    .Y(_04134_)
  );
  sg13g2_nor2_1 _14235_ (
    .A(_01187_),
    .B(_04134_),
    .Y(_04135_)
  );
  sg13g2_o21ai_1 _14236_ (
    .A1(_03842_),
    .A2(_00559_),
    .B1(addr_i_3_),
    .Y(_04136_)
  );
  sg13g2_nand4_1 _14237_ (
    .A(addr_i_7_),
    .B(_00831_),
    .C(_01425_),
    .D(_04136_),
    .Y(_04137_)
  );
  sg13g2_nand3_1 _14238_ (
    .A(_05811_),
    .B(_04041_),
    .C(_01462_),
    .Y(_04138_)
  );
  sg13g2_nor2_1 _14239_ (
    .A(_07757_),
    .B(_09393_),
    .Y(_04139_)
  );
  sg13g2_nand2_1 _14240_ (
    .A(_00744_),
    .B(_00985_),
    .Y(_04141_)
  );
  sg13g2_a21oi_1 _14241_ (
    .A1(_06088_),
    .A2(_04141_),
    .B1(addr_i_3_),
    .Y(_04142_)
  );
  sg13g2_a221oi_1 _14242_ (
    .A1(_04137_),
    .A2(_04138_),
    .B1(_04139_),
    .B2(addr_i_3_),
    .C1(_04142_),
    .Y(_04143_)
  );
  sg13g2_a22oi_1 _14243_ (
    .A1(_00402_),
    .A2(_04135_),
    .B1(_04143_),
    .B2(addr_i_8_),
    .Y(_04144_)
  );
  sg13g2_nand2_1 _14244_ (
    .A(_07812_),
    .B(_05689_),
    .Y(_04145_)
  );
  sg13g2_o21ai_1 _14245_ (
    .A1(addr_i_2_),
    .A2(_01019_),
    .B1(_04145_),
    .Y(_04146_)
  );
  sg13g2_nand2_1 _14246_ (
    .A(addr_i_8_),
    .B(_01543_),
    .Y(_04147_)
  );
  sg13g2_nor2_1 _14247_ (
    .A(_05535_),
    .B(_00405_),
    .Y(_04148_)
  );
  sg13g2_a22oi_1 _14248_ (
    .A1(_09474_),
    .A2(_04146_),
    .B1(_04147_),
    .B2(_04148_),
    .Y(_04149_)
  );
  sg13g2_or3_1 _14249_ (
    .A(addr_i_9_),
    .B(_04144_),
    .C(_04149_),
    .X(_04150_)
  );
  sg13g2_nor2_1 _14250_ (
    .A(_00497_),
    .B(_01666_),
    .Y(_04152_)
  );
  sg13g2_o21ai_1 _14251_ (
    .A1(_04152_),
    .A2(_01360_),
    .B1(addr_i_9_),
    .Y(_04153_)
  );
  sg13g2_a21oi_1 _14252_ (
    .A1(_04150_),
    .A2(_04153_),
    .B1(addr_i_10_),
    .Y(_04154_)
  );
  sg13g2_o21ai_1 _14253_ (
    .A1(_04133_),
    .A2(_04154_),
    .B1(addr_i_12_),
    .Y(_04155_)
  );
  sg13g2_nand2_1 _14254_ (
    .A(_01279_),
    .B(_00853_),
    .Y(_04156_)
  );
  sg13g2_nor3_1 _14255_ (
    .A(addr_i_3_),
    .B(_00491_),
    .C(_01216_),
    .Y(_04157_)
  );
  sg13g2_nor2_1 _14256_ (
    .A(_02179_),
    .B(_04157_),
    .Y(_04158_)
  );
  sg13g2_a21oi_1 _14257_ (
    .A1(_04156_),
    .A2(_04158_),
    .B1(addr_i_9_),
    .Y(_04159_)
  );
  sg13g2_o21ai_1 _14258_ (
    .A1(_00115_),
    .A2(_02560_),
    .B1(_02497_),
    .Y(_04160_)
  );
  sg13g2_a21oi_1 _14259_ (
    .A1(_00762_),
    .A2(_09478_),
    .B1(_03652_),
    .Y(_04161_)
  );
  sg13g2_a21oi_1 _14260_ (
    .A1(addr_i_7_),
    .A2(_04160_),
    .B1(_04161_),
    .Y(_04163_)
  );
  sg13g2_o21ai_1 _14261_ (
    .A1(addr_i_2_),
    .A2(_00000_),
    .B1(addr_i_4_),
    .Y(_04164_)
  );
  sg13g2_a21oi_1 _14262_ (
    .A1(_01267_),
    .A2(_04164_),
    .B1(addr_i_3_),
    .Y(_04165_)
  );
  sg13g2_o21ai_1 _14263_ (
    .A1(_05258_),
    .A2(_03632_),
    .B1(addr_i_3_),
    .Y(_04166_)
  );
  sg13g2_nand2_1 _14264_ (
    .A(_09260_),
    .B(_04166_),
    .Y(_04167_)
  );
  sg13g2_o21ai_1 _14265_ (
    .A1(_04165_),
    .A2(_04167_),
    .B1(_01475_),
    .Y(_04168_)
  );
  sg13g2_o21ai_1 _14266_ (
    .A1(addr_i_6_),
    .A2(_04163_),
    .B1(_04168_),
    .Y(_04169_)
  );
  sg13g2_nand2_1 _14267_ (
    .A(_00626_),
    .B(_02103_),
    .Y(_04170_)
  );
  sg13g2_a22oi_1 _14268_ (
    .A1(addr_i_3_),
    .A2(_02278_),
    .B1(_00885_),
    .B2(_08299_),
    .Y(_04171_)
  );
  sg13g2_o21ai_1 _14269_ (
    .A1(addr_i_7_),
    .A2(_04171_),
    .B1(_03575_),
    .Y(_04172_)
  );
  sg13g2_nand2_1 _14270_ (
    .A(_01794_),
    .B(_04172_),
    .Y(_04175_)
  );
  sg13g2_a21oi_1 _14271_ (
    .A1(_08376_),
    .A2(_00049_),
    .B1(_02459_),
    .Y(_04176_)
  );
  sg13g2_o21ai_1 _14272_ (
    .A1(_01514_),
    .A2(_01673_),
    .B1(_01152_),
    .Y(_04177_)
  );
  sg13g2_o21ai_1 _14273_ (
    .A1(_04176_),
    .A2(_04177_),
    .B1(addr_i_4_),
    .Y(_04178_)
  );
  sg13g2_nand4_1 _14274_ (
    .A(addr_i_8_),
    .B(_04170_),
    .C(_04175_),
    .D(_04178_),
    .Y(_04179_)
  );
  sg13g2_o21ai_1 _14275_ (
    .A1(addr_i_8_),
    .A2(_04169_),
    .B1(_04179_),
    .Y(_04180_)
  );
  sg13g2_nor2_1 _14276_ (
    .A(_00967_),
    .B(_00939_),
    .Y(_04181_)
  );
  sg13g2_a22oi_1 _14277_ (
    .A1(_01520_),
    .A2(_00473_),
    .B1(_04181_),
    .B2(_03260_),
    .Y(_04182_)
  );
  sg13g2_a22oi_1 _14278_ (
    .A1(addr_i_4_),
    .A2(_07480_),
    .B1(_01387_),
    .B2(addr_i_3_),
    .Y(_04183_)
  );
  sg13g2_o21ai_1 _14279_ (
    .A1(_04182_),
    .A2(_04183_),
    .B1(_02467_),
    .Y(_04184_)
  );
  sg13g2_nand2_1 _14280_ (
    .A(addr_i_4_),
    .B(_01373_),
    .Y(_04186_)
  );
  sg13g2_nand2_1 _14281_ (
    .A(_02118_),
    .B(_00358_),
    .Y(_04187_)
  );
  sg13g2_o21ai_1 _14282_ (
    .A1(_04186_),
    .A2(_03012_),
    .B1(_04187_),
    .Y(_04188_)
  );
  sg13g2_o21ai_1 _14283_ (
    .A1(_01034_),
    .A2(_04188_),
    .B1(addr_i_9_),
    .Y(_04189_)
  );
  sg13g2_a21oi_1 _14284_ (
    .A1(addr_i_6_),
    .A2(_00719_),
    .B1(_08155_),
    .Y(_04190_)
  );
  sg13g2_buf_1 _14285_ (
    .A(_03919_),
    .X(_04191_)
  );
  sg13g2_o21ai_1 _14286_ (
    .A1(_00561_),
    .A2(_04190_),
    .B1(_04191_),
    .Y(_04192_)
  );
  sg13g2_a22oi_1 _14287_ (
    .A1(_00999_),
    .A2(_01808_),
    .B1(_01819_),
    .B2(_01285_),
    .Y(_04193_)
  );
  sg13g2_nand2_1 _14288_ (
    .A(_04192_),
    .B(_04193_),
    .Y(_04194_)
  );
  sg13g2_nand2b_1 _14289_ (
    .A_N(_03905_),
    .B(addr_i_3_),
    .Y(_04195_)
  );
  sg13g2_o21ai_1 _14290_ (
    .A1(_00491_),
    .A2(_01896_),
    .B1(addr_i_6_),
    .Y(_04197_)
  );
  sg13g2_a21oi_1 _14291_ (
    .A1(_04195_),
    .A2(_04197_),
    .B1(addr_i_4_),
    .Y(_04198_)
  );
  sg13g2_a22oi_1 _14292_ (
    .A1(_00360_),
    .A2(_00917_),
    .B1(_01402_),
    .B2(addr_i_3_),
    .Y(_04199_)
  );
  sg13g2_o21ai_1 _14293_ (
    .A1(addr_i_5_),
    .A2(_01014_),
    .B1(addr_i_4_),
    .Y(_04200_)
  );
  sg13g2_a22oi_1 _14294_ (
    .A1(addr_i_2_),
    .A2(_06132_),
    .B1(_06398_),
    .B2(_06419_),
    .Y(_04201_)
  );
  sg13g2_and2_1 _14295_ (
    .A(_04200_),
    .B(_04201_),
    .X(_04202_)
  );
  sg13g2_o21ai_1 _14296_ (
    .A1(_04199_),
    .A2(_04202_),
    .B1(_01861_),
    .Y(_04203_)
  );
  sg13g2_o21ai_1 _14297_ (
    .A1(_04194_),
    .A2(_04198_),
    .B1(_04203_),
    .Y(_04204_)
  );
  sg13g2_a22oi_1 _14298_ (
    .A1(_00277_),
    .A2(_04184_),
    .B1(_04189_),
    .B2(_04204_),
    .Y(_04205_)
  );
  sg13g2_a22oi_1 _14299_ (
    .A1(_04159_),
    .A2(_04180_),
    .B1(_04205_),
    .B2(addr_i_10_),
    .Y(_04206_)
  );
  sg13g2_nand2_1 _14300_ (
    .A(addr_i_2_),
    .B(_02405_),
    .Y(_04208_)
  );
  sg13g2_o21ai_1 _14301_ (
    .A1(_01212_),
    .A2(_01616_),
    .B1(_04208_),
    .Y(_04209_)
  );
  sg13g2_o21ai_1 _14302_ (
    .A1(_01231_),
    .A2(_01232_),
    .B1(_00261_),
    .Y(_04210_)
  );
  sg13g2_a21oi_1 _14303_ (
    .A1(_03575_),
    .A2(_04210_),
    .B1(addr_i_3_),
    .Y(_04211_)
  );
  sg13g2_a22oi_1 _14304_ (
    .A1(addr_i_3_),
    .A2(_04209_),
    .B1(_04211_),
    .B2(_00977_),
    .Y(_04212_)
  );
  sg13g2_nand2_1 _14305_ (
    .A(_00434_),
    .B(_00620_),
    .Y(_04213_)
  );
  sg13g2_nand2_1 _14306_ (
    .A(_00453_),
    .B(_01337_),
    .Y(_04214_)
  );
  sg13g2_a21oi_1 _14307_ (
    .A1(_08221_),
    .A2(_02089_),
    .B1(addr_i_3_),
    .Y(_04215_)
  );
  sg13g2_a221oi_1 _14308_ (
    .A1(addr_i_5_),
    .A2(_04213_),
    .B1(_04214_),
    .B2(addr_i_3_),
    .C1(_04215_),
    .Y(_04216_)
  );
  sg13g2_mux2_1 _14309_ (
    .A0(_04212_),
    .A1(_04216_),
    .S(addr_i_4_),
    .X(_04217_)
  );
  sg13g2_nor2_1 _14310_ (
    .A(_01262_),
    .B(_00080_),
    .Y(_04219_)
  );
  sg13g2_o21ai_1 _14311_ (
    .A1(_00247_),
    .A2(_04219_),
    .B1(_03260_),
    .Y(_04220_)
  );
  sg13g2_nand3_1 _14312_ (
    .A(_00186_),
    .B(_03778_),
    .C(_04220_),
    .Y(_04221_)
  );
  sg13g2_nand2_1 _14313_ (
    .A(_07812_),
    .B(_00008_),
    .Y(_04222_)
  );
  sg13g2_nand2_1 _14314_ (
    .A(_00844_),
    .B(_01580_),
    .Y(_04223_)
  );
  sg13g2_a21oi_1 _14315_ (
    .A1(_04222_),
    .A2(_04223_),
    .B1(addr_i_6_),
    .Y(_04224_)
  );
  sg13g2_a21oi_1 _14316_ (
    .A1(_03446_),
    .A2(_01066_),
    .B1(addr_i_4_),
    .Y(_04225_)
  );
  sg13g2_a221oi_1 _14317_ (
    .A1(_01227_),
    .A2(_03905_),
    .B1(_04225_),
    .B2(_02530_),
    .C1(_00945_),
    .Y(_04226_)
  );
  sg13g2_a21oi_1 _14318_ (
    .A1(_00073_),
    .A2(_06276_),
    .B1(_00782_),
    .Y(_04227_)
  );
  sg13g2_o21ai_1 _14319_ (
    .A1(addr_i_7_),
    .A2(_04226_),
    .B1(_04227_),
    .Y(_04228_)
  );
  sg13g2_a22oi_1 _14320_ (
    .A1(addr_i_6_),
    .A2(_04221_),
    .B1(_04224_),
    .B2(_04228_),
    .Y(_04230_)
  );
  sg13g2_a22oi_1 _14321_ (
    .A1(_00114_),
    .A2(_04217_),
    .B1(_04230_),
    .B2(_00109_),
    .Y(_04231_)
  );
  sg13g2_o21ai_1 _14322_ (
    .A1(addr_i_3_),
    .A2(_01212_),
    .B1(_04207_),
    .Y(_04232_)
  );
  sg13g2_a21oi_1 _14323_ (
    .A1(_04296_),
    .A2(_03424_),
    .B1(_01514_),
    .Y(_04233_)
  );
  sg13g2_a21o_1 _14324_ (
    .A1(addr_i_6_),
    .A2(_04232_),
    .B1(_04233_),
    .X(_04234_)
  );
  sg13g2_o21ai_1 _14325_ (
    .A1(_06950_),
    .A2(_05645_),
    .B1(addr_i_3_),
    .Y(_04235_)
  );
  sg13g2_nand2_1 _14326_ (
    .A(_00190_),
    .B(_02080_),
    .Y(_04236_)
  );
  sg13g2_nand3_1 _14327_ (
    .A(_01224_),
    .B(_04235_),
    .C(_04236_),
    .Y(_04237_)
  );
  sg13g2_nor2_1 _14328_ (
    .A(_01972_),
    .B(_02848_),
    .Y(_04238_)
  );
  sg13g2_nor2_1 _14329_ (
    .A(_00878_),
    .B(_04238_),
    .Y(_04239_)
  );
  sg13g2_a221oi_1 _14330_ (
    .A1(addr_i_4_),
    .A2(_04234_),
    .B1(_04237_),
    .B2(addr_i_2_),
    .C1(_04239_),
    .Y(_04241_)
  );
  sg13g2_o21ai_1 _14331_ (
    .A1(_02040_),
    .A2(_04241_),
    .B1(_01640_),
    .Y(_04242_)
  );
  sg13g2_o21ai_1 _14332_ (
    .A1(_06010_),
    .A2(_09499_),
    .B1(addr_i_2_),
    .Y(_04243_)
  );
  sg13g2_o21ai_1 _14333_ (
    .A1(addr_i_7_),
    .A2(_00666_),
    .B1(_01441_),
    .Y(_04244_)
  );
  sg13g2_nand2_1 _14334_ (
    .A(_01630_),
    .B(_04244_),
    .Y(_04245_)
  );
  sg13g2_nor2_1 _14335_ (
    .A(_03809_),
    .B(_02152_),
    .Y(_04246_)
  );
  sg13g2_o21ai_1 _14336_ (
    .A1(_07425_),
    .A2(_04246_),
    .B1(addr_i_4_),
    .Y(_04247_)
  );
  sg13g2_nand3_1 _14337_ (
    .A(_04243_),
    .B(_04245_),
    .C(_04247_),
    .Y(_04248_)
  );
  sg13g2_nand2_1 _14338_ (
    .A(_00403_),
    .B(_00573_),
    .Y(_04249_)
  );
  sg13g2_a22oi_1 _14339_ (
    .A1(addr_i_7_),
    .A2(_04249_),
    .B1(_03572_),
    .B2(_00068_),
    .Y(_04250_)
  );
  sg13g2_nand2_1 _14340_ (
    .A(addr_i_4_),
    .B(_03110_),
    .Y(_04252_)
  );
  sg13g2_a21oi_1 _14341_ (
    .A1(_03226_),
    .A2(_04252_),
    .B1(addr_i_7_),
    .Y(_04253_)
  );
  sg13g2_a22oi_1 _14342_ (
    .A1(_00386_),
    .A2(_00128_),
    .B1(_04253_),
    .B2(addr_i_2_),
    .Y(_04254_)
  );
  sg13g2_nor3_1 _14343_ (
    .A(addr_i_3_),
    .B(_04250_),
    .C(_04254_),
    .Y(_04255_)
  );
  sg13g2_a21oi_1 _14344_ (
    .A1(addr_i_3_),
    .A2(_04248_),
    .B1(_04255_),
    .Y(_04256_)
  );
  sg13g2_nor2_1 _14345_ (
    .A(_04036_),
    .B(_04256_),
    .Y(_04257_)
  );
  sg13g2_nor4_1 _14346_ (
    .A(_04206_),
    .B(_04231_),
    .C(_04242_),
    .D(_04257_),
    .Y(_04258_)
  );
  sg13g2_a21oi_1 _14347_ (
    .A1(_02404_),
    .A2(_05501_),
    .B1(_00156_),
    .Y(_04259_)
  );
  sg13g2_o21ai_1 _14348_ (
    .A1(addr_i_5_),
    .A2(_04259_),
    .B1(_00443_),
    .Y(_04260_)
  );
  sg13g2_a21oi_1 _14349_ (
    .A1(addr_i_4_),
    .A2(_00581_),
    .B1(addr_i_3_),
    .Y(_04261_)
  );
  sg13g2_o21ai_1 _14350_ (
    .A1(_00268_),
    .A2(_04261_),
    .B1(_02501_),
    .Y(_04263_)
  );
  sg13g2_nand2_1 _14351_ (
    .A(addr_i_9_),
    .B(_04263_),
    .Y(_04264_)
  );
  sg13g2_a21oi_1 _14352_ (
    .A1(_07469_),
    .A2(_00725_),
    .B1(_09038_),
    .Y(_04265_)
  );
  sg13g2_o21ai_1 _14353_ (
    .A1(_00587_),
    .A2(_04265_),
    .B1(addr_i_4_),
    .Y(_04266_)
  );
  sg13g2_a21oi_1 _14354_ (
    .A1(_00739_),
    .A2(_04266_),
    .B1(_07403_),
    .Y(_04267_)
  );
  sg13g2_a22oi_1 _14355_ (
    .A1(_02498_),
    .A2(_04260_),
    .B1(_04264_),
    .B2(_04267_),
    .Y(_04268_)
  );
  sg13g2_a21oi_1 _14356_ (
    .A1(_03798_),
    .A2(_00462_),
    .B1(addr_i_3_),
    .Y(_04269_)
  );
  sg13g2_o21ai_1 _14357_ (
    .A1(_06972_),
    .A2(_00813_),
    .B1(_03413_),
    .Y(_04270_)
  );
  sg13g2_o21ai_1 _14358_ (
    .A1(_04269_),
    .A2(_04270_),
    .B1(addr_i_4_),
    .Y(_04271_)
  );
  sg13g2_o21ai_1 _14359_ (
    .A1(_01153_),
    .A2(_03589_),
    .B1(addr_i_3_),
    .Y(_04272_)
  );
  sg13g2_nand3_1 _14360_ (
    .A(_02810_),
    .B(_04271_),
    .C(_04272_),
    .Y(_04274_)
  );
  sg13g2_a21oi_1 _14361_ (
    .A1(_02471_),
    .A2(_01203_),
    .B1(_02001_),
    .Y(_04275_)
  );
  sg13g2_nor2_1 _14362_ (
    .A(_03776_),
    .B(_09509_),
    .Y(_04276_)
  );
  sg13g2_a22oi_1 _14363_ (
    .A1(addr_i_6_),
    .A2(_04274_),
    .B1(_04275_),
    .B2(_04276_),
    .Y(_04277_)
  );
  sg13g2_or2_1 _14364_ (
    .A(addr_i_8_),
    .B(_04277_),
    .X(_04278_)
  );
  sg13g2_nor3_1 _14365_ (
    .A(_04949_),
    .B(_09502_),
    .C(_00721_),
    .Y(_04279_)
  );
  sg13g2_o21ai_1 _14366_ (
    .A1(_01065_),
    .A2(_01754_),
    .B1(_04279_),
    .Y(_04280_)
  );
  sg13g2_nor2_1 _14367_ (
    .A(_04418_),
    .B(_00964_),
    .Y(_04281_)
  );
  sg13g2_nand2_1 _14368_ (
    .A(_07326_),
    .B(_04429_),
    .Y(_04282_)
  );
  sg13g2_nor4_1 _14369_ (
    .A(_00205_),
    .B(_04281_),
    .C(_02055_),
    .D(_04282_),
    .Y(_04283_)
  );
  sg13g2_nor2_1 _14370_ (
    .A(addr_i_3_),
    .B(_04283_),
    .Y(_04286_)
  );
  sg13g2_a22oi_1 _14371_ (
    .A1(addr_i_3_),
    .A2(_04280_),
    .B1(_04286_),
    .B2(_02794_),
    .Y(_04287_)
  );
  sg13g2_or2_1 _14372_ (
    .A(_05734_),
    .B(_01337_),
    .X(_04288_)
  );
  sg13g2_o21ai_1 _14373_ (
    .A1(_03676_),
    .A2(_02503_),
    .B1(_00099_),
    .Y(_04289_)
  );
  sg13g2_nand4_1 _14374_ (
    .A(_03687_),
    .B(_03707_),
    .C(_04288_),
    .D(_04289_),
    .Y(_04290_)
  );
  sg13g2_nand2_1 _14375_ (
    .A(_08796_),
    .B(_08852_),
    .Y(_04291_)
  );
  sg13g2_nand2_1 _14376_ (
    .A(_00086_),
    .B(_03110_),
    .Y(_04292_)
  );
  sg13g2_o21ai_1 _14377_ (
    .A1(addr_i_2_),
    .A2(_03172_),
    .B1(_02369_),
    .Y(_04293_)
  );
  sg13g2_nand3_1 _14378_ (
    .A(_04291_),
    .B(_04292_),
    .C(_04293_),
    .Y(_04294_)
  );
  sg13g2_nand2_1 _14379_ (
    .A(_04926_),
    .B(_04860_),
    .Y(_04295_)
  );
  sg13g2_a21oi_1 _14380_ (
    .A1(_01543_),
    .A2(_04295_),
    .B1(_00522_),
    .Y(_04297_)
  );
  sg13g2_a221oi_1 _14381_ (
    .A1(_02287_),
    .A2(_04290_),
    .B1(_04294_),
    .B2(addr_i_4_),
    .C1(_04297_),
    .Y(_04298_)
  );
  sg13g2_nor2_1 _14382_ (
    .A(addr_i_8_),
    .B(_04298_),
    .Y(_04299_)
  );
  sg13g2_a22oi_1 _14383_ (
    .A1(addr_i_8_),
    .A2(_04287_),
    .B1(_04299_),
    .B2(addr_i_9_),
    .Y(_04300_)
  );
  sg13g2_a22oi_1 _14384_ (
    .A1(_04268_),
    .A2(_04278_),
    .B1(addr_i_10_),
    .B2(_04300_),
    .Y(_04301_)
  );
  sg13g2_o21ai_1 _14385_ (
    .A1(_03540_),
    .A2(_00557_),
    .B1(_00915_),
    .Y(_04302_)
  );
  sg13g2_a22oi_1 _14386_ (
    .A1(_02105_),
    .A2(_04302_),
    .B1(_02873_),
    .B2(addr_i_4_),
    .Y(_04303_)
  );
  sg13g2_o21ai_1 _14387_ (
    .A1(_00158_),
    .A2(_02218_),
    .B1(_08254_),
    .Y(_04304_)
  );
  sg13g2_a22oi_1 _14388_ (
    .A1(addr_i_7_),
    .A2(_04304_),
    .B1(_01837_),
    .B2(_01131_),
    .Y(_04305_)
  );
  sg13g2_a21oi_1 _14389_ (
    .A1(_00016_),
    .A2(_04628_),
    .B1(addr_i_3_),
    .Y(_04306_)
  );
  sg13g2_a22oi_1 _14390_ (
    .A1(_00442_),
    .A2(_02382_),
    .B1(_04306_),
    .B2(_06950_),
    .Y(_04308_)
  );
  sg13g2_nand2b_1 _14391_ (
    .A_N(_04308_),
    .B(addr_i_6_),
    .Y(_04309_)
  );
  sg13g2_o21ai_1 _14392_ (
    .A1(_04303_),
    .A2(_04305_),
    .B1(_04309_),
    .Y(_04310_)
  );
  sg13g2_o21ai_1 _14393_ (
    .A1(_01107_),
    .A2(_03112_),
    .B1(addr_i_7_),
    .Y(_04311_)
  );
  sg13g2_a21oi_1 _14394_ (
    .A1(_04384_),
    .A2(_01273_),
    .B1(addr_i_4_),
    .Y(_04312_)
  );
  sg13g2_nor2_1 _14395_ (
    .A(_00046_),
    .B(_04312_),
    .Y(_04313_)
  );
  sg13g2_nor4_1 _14396_ (
    .A(addr_i_3_),
    .B(_06751_),
    .C(_01567_),
    .D(_01732_),
    .Y(_04314_)
  );
  sg13g2_a21oi_1 _14397_ (
    .A1(_04311_),
    .A2(_04313_),
    .B1(_04314_),
    .Y(_04315_)
  );
  sg13g2_nor2_1 _14398_ (
    .A(_05845_),
    .B(_02558_),
    .Y(_04316_)
  );
  sg13g2_a21oi_1 _14399_ (
    .A1(_00700_),
    .A2(_00384_),
    .B1(_04316_),
    .Y(_04317_)
  );
  sg13g2_o21ai_1 _14400_ (
    .A1(_01747_),
    .A2(_03742_),
    .B1(addr_i_4_),
    .Y(_04319_)
  );
  sg13g2_o21ai_1 _14401_ (
    .A1(_00840_),
    .A2(_04317_),
    .B1(_04319_),
    .Y(_04320_)
  );
  sg13g2_nor3_1 _14402_ (
    .A(addr_i_8_),
    .B(_04315_),
    .C(_04320_),
    .Y(_04321_)
  );
  sg13g2_a22oi_1 _14403_ (
    .A1(addr_i_8_),
    .A2(_04310_),
    .B1(_04321_),
    .B2(_04705_),
    .Y(_04322_)
  );
  sg13g2_nor4_1 _14404_ (
    .A(_00977_),
    .B(_00238_),
    .C(_05634_),
    .D(_02983_),
    .Y(_04323_)
  );
  sg13g2_a21oi_1 _14405_ (
    .A1(_01273_),
    .A2(_01441_),
    .B1(_00059_),
    .Y(_04324_)
  );
  sg13g2_nor2_1 _14406_ (
    .A(_04215_),
    .B(_04324_),
    .Y(_04325_)
  );
  sg13g2_o21ai_1 _14407_ (
    .A1(addr_i_4_),
    .A2(_04323_),
    .B1(_04325_),
    .Y(_04326_)
  );
  sg13g2_nor3_1 _14408_ (
    .A(_03617_),
    .B(_00023_),
    .C(_04326_),
    .Y(_04327_)
  );
  sg13g2_nand2_1 _14409_ (
    .A(_03798_),
    .B(_01757_),
    .Y(_04328_)
  );
  sg13g2_nand2_1 _14410_ (
    .A(addr_i_3_),
    .B(_04328_),
    .Y(_04330_)
  );
  sg13g2_nand3_1 _14411_ (
    .A(_00910_),
    .B(_01070_),
    .C(_03575_),
    .Y(_04331_)
  );
  sg13g2_nand3_1 _14412_ (
    .A(addr_i_4_),
    .B(_04330_),
    .C(_04331_),
    .Y(_04332_)
  );
  sg13g2_nand2_1 _14413_ (
    .A(addr_i_2_),
    .B(_00025_),
    .Y(_04333_)
  );
  sg13g2_a22oi_1 _14414_ (
    .A1(_08696_),
    .A2(_04333_),
    .B1(_00096_),
    .B2(_00059_),
    .Y(_04334_)
  );
  sg13g2_nor3_1 _14415_ (
    .A(addr_i_3_),
    .B(addr_i_5_),
    .C(_01507_),
    .Y(_04335_)
  );
  sg13g2_nand2_1 _14416_ (
    .A(addr_i_6_),
    .B(_02618_),
    .Y(_04336_)
  );
  sg13g2_o21ai_1 _14417_ (
    .A1(_04334_),
    .A2(_04335_),
    .B1(_04336_),
    .Y(_04337_)
  );
  sg13g2_a21oi_1 _14418_ (
    .A1(_01175_),
    .A2(_02149_),
    .B1(_06419_),
    .Y(_04338_)
  );
  sg13g2_a22oi_1 _14419_ (
    .A1(_01972_),
    .A2(_08774_),
    .B1(_04338_),
    .B2(addr_i_4_),
    .Y(_04339_)
  );
  sg13g2_a21oi_1 _14420_ (
    .A1(_04396_),
    .A2(_00687_),
    .B1(_00293_),
    .Y(_04341_)
  );
  sg13g2_o21ai_1 _14421_ (
    .A1(_01159_),
    .A2(_04341_),
    .B1(_00799_),
    .Y(_04342_)
  );
  sg13g2_a221oi_1 _14422_ (
    .A1(addr_i_4_),
    .A2(_04337_),
    .B1(_04339_),
    .B2(_04342_),
    .C1(addr_i_8_),
    .Y(_04343_)
  );
  sg13g2_a22oi_1 _14423_ (
    .A1(_04327_),
    .A2(_04332_),
    .B1(addr_i_9_),
    .B2(_04343_),
    .Y(_04344_)
  );
  sg13g2_nor3_1 _14424_ (
    .A(_01773_),
    .B(_04322_),
    .C(_04344_),
    .Y(_04345_)
  );
  sg13g2_nor3_1 _14425_ (
    .A(_03040_),
    .B(_04301_),
    .C(_04345_),
    .Y(_04346_)
  );
  sg13g2_a21oi_1 _14426_ (
    .A1(_00370_),
    .A2(_00125_),
    .B1(_08852_),
    .Y(_04347_)
  );
  sg13g2_o21ai_1 _14427_ (
    .A1(_02801_),
    .A2(_04347_),
    .B1(_04650_),
    .Y(_04348_)
  );
  sg13g2_a21oi_1 _14428_ (
    .A1(_05745_),
    .A2(_00014_),
    .B1(_01663_),
    .Y(_04349_)
  );
  sg13g2_o21ai_1 _14429_ (
    .A1(_00731_),
    .A2(_00972_),
    .B1(_04349_),
    .Y(_04350_)
  );
  sg13g2_o21ai_1 _14430_ (
    .A1(addr_i_6_),
    .A2(_07237_),
    .B1(_00064_),
    .Y(_04352_)
  );
  sg13g2_nand3_1 _14431_ (
    .A(addr_i_4_),
    .B(_03765_),
    .C(_01055_),
    .Y(_04353_)
  );
  sg13g2_nand4_1 _14432_ (
    .A(_00535_),
    .B(_01406_),
    .C(_04352_),
    .D(_04353_),
    .Y(_04354_)
  );
  sg13g2_nand2_1 _14433_ (
    .A(addr_i_2_),
    .B(_02591_),
    .Y(_04355_)
  );
  sg13g2_nand3_1 _14434_ (
    .A(addr_i_3_),
    .B(_01175_),
    .C(_04355_),
    .Y(_04356_)
  );
  sg13g2_a21o_1 _14435_ (
    .A1(_04354_),
    .A2(_04356_),
    .B1(_01274_),
    .X(_04357_)
  );
  sg13g2_and4_1 _14436_ (
    .A(_00374_),
    .B(_04348_),
    .C(_04350_),
    .D(_04357_),
    .X(_04358_)
  );
  sg13g2_nand3_1 _14437_ (
    .A(addr_i_3_),
    .B(_04063_),
    .C(_00148_),
    .Y(_04359_)
  );
  sg13g2_a21oi_1 _14438_ (
    .A1(_01397_),
    .A2(_04359_),
    .B1(_02344_),
    .Y(_04360_)
  );
  sg13g2_nor3_1 _14439_ (
    .A(addr_i_6_),
    .B(_02297_),
    .C(_01571_),
    .Y(_04361_)
  );
  sg13g2_o21ai_1 _14440_ (
    .A1(_04360_),
    .A2(_04361_),
    .B1(_01666_),
    .Y(_04363_)
  );
  sg13g2_a21o_1 _14441_ (
    .A1(_01073_),
    .A2(_04077_),
    .B1(addr_i_2_),
    .X(_04364_)
  );
  sg13g2_a22oi_1 _14442_ (
    .A1(addr_i_4_),
    .A2(_09448_),
    .B1(_01957_),
    .B2(_00860_),
    .Y(_04365_)
  );
  sg13g2_o21ai_1 _14443_ (
    .A1(addr_i_3_),
    .A2(_01094_),
    .B1(_01432_),
    .Y(_04366_)
  );
  sg13g2_nand2_1 _14444_ (
    .A(_00915_),
    .B(_00333_),
    .Y(_04367_)
  );
  sg13g2_a221oi_1 _14445_ (
    .A1(addr_i_4_),
    .A2(_04366_),
    .B1(_04367_),
    .B2(_01215_),
    .C1(_06276_),
    .Y(_04368_)
  );
  sg13g2_nor2_1 _14446_ (
    .A(_03227_),
    .B(_04368_),
    .Y(_04369_)
  );
  sg13g2_a22oi_1 _14447_ (
    .A1(_04364_),
    .A2(_04365_),
    .B1(_09315_),
    .B2(_04369_),
    .Y(_04370_)
  );
  sg13g2_nand2_1 _14448_ (
    .A(_00637_),
    .B(_08763_),
    .Y(_04371_)
  );
  sg13g2_nand3_1 _14449_ (
    .A(_09415_),
    .B(_01912_),
    .C(_04371_),
    .Y(_04372_)
  );
  sg13g2_a21oi_1 _14450_ (
    .A1(_01729_),
    .A2(_02683_),
    .B1(addr_i_3_),
    .Y(_04374_)
  );
  sg13g2_a22oi_1 _14451_ (
    .A1(addr_i_3_),
    .A2(_04372_),
    .B1(_04374_),
    .B2(_00206_),
    .Y(_04375_)
  );
  sg13g2_nor2_1 _14452_ (
    .A(_01099_),
    .B(_04375_),
    .Y(_04376_)
  );
  sg13g2_nor3_1 _14453_ (
    .A(_00024_),
    .B(_00616_),
    .C(_01281_),
    .Y(_04377_)
  );
  sg13g2_o21ai_1 _14454_ (
    .A1(_01014_),
    .A2(_02443_),
    .B1(_08741_),
    .Y(_04378_)
  );
  sg13g2_o21ai_1 _14455_ (
    .A1(_02441_),
    .A2(_03566_),
    .B1(addr_i_3_),
    .Y(_04379_)
  );
  sg13g2_a21oi_1 _14456_ (
    .A1(_04378_),
    .A2(_04379_),
    .B1(_00445_),
    .Y(_04380_)
  );
  sg13g2_o21ai_1 _14457_ (
    .A1(_04377_),
    .A2(_04380_),
    .B1(_01118_),
    .Y(_04381_)
  );
  sg13g2_nor2b_1 _14458_ (
    .A(_04376_),
    .B_N(_04381_),
    .Y(_04382_)
  );
  sg13g2_a221oi_1 _14459_ (
    .A1(_04358_),
    .A2(_04363_),
    .B1(_04370_),
    .B2(_04382_),
    .C1(addr_i_10_),
    .Y(_04383_)
  );
  sg13g2_o21ai_1 _14460_ (
    .A1(addr_i_2_),
    .A2(_09485_),
    .B1(_00915_),
    .Y(_04385_)
  );
  sg13g2_a21oi_1 _14461_ (
    .A1(_00965_),
    .A2(_08520_),
    .B1(_00260_),
    .Y(_04386_)
  );
  sg13g2_a22oi_1 _14462_ (
    .A1(_05402_),
    .A2(_04385_),
    .B1(_04386_),
    .B2(_01587_),
    .Y(_04387_)
  );
  sg13g2_a21oi_1 _14463_ (
    .A1(_00586_),
    .A2(_03413_),
    .B1(_01120_),
    .Y(_04388_)
  );
  sg13g2_a21oi_1 _14464_ (
    .A1(_01603_),
    .A2(_01834_),
    .B1(_05856_),
    .Y(_04389_)
  );
  sg13g2_o21ai_1 _14465_ (
    .A1(_04388_),
    .A2(_04389_),
    .B1(addr_i_6_),
    .Y(_04390_)
  );
  sg13g2_o21ai_1 _14466_ (
    .A1(addr_i_3_),
    .A2(_04387_),
    .B1(_04390_),
    .Y(_04391_)
  );
  sg13g2_o21ai_1 _14467_ (
    .A1(_00015_),
    .A2(_02873_),
    .B1(_02277_),
    .Y(_04392_)
  );
  sg13g2_nand3b_1 _14468_ (
    .A_N(_04391_),
    .B(_04392_),
    .C(_01601_),
    .Y(_04393_)
  );
  sg13g2_a21oi_1 _14469_ (
    .A1(_09476_),
    .A2(_00453_),
    .B1(addr_i_3_),
    .Y(_04394_)
  );
  sg13g2_o21ai_1 _14470_ (
    .A1(_00850_),
    .A2(_04394_),
    .B1(_02257_),
    .Y(_04397_)
  );
  sg13g2_o21ai_1 _14471_ (
    .A1(_00959_),
    .A2(_02652_),
    .B1(addr_i_5_),
    .Y(_04398_)
  );
  sg13g2_nor2_1 _14472_ (
    .A(addr_i_7_),
    .B(_07658_),
    .Y(_04399_)
  );
  sg13g2_nor2_1 _14473_ (
    .A(_07160_),
    .B(_02459_),
    .Y(_04400_)
  );
  sg13g2_a21oi_1 _14474_ (
    .A1(_01653_),
    .A2(_04399_),
    .B1(_04400_),
    .Y(_04401_)
  );
  sg13g2_nand2_1 _14475_ (
    .A(_04398_),
    .B(_04401_),
    .Y(_04402_)
  );
  sg13g2_nor3_1 _14476_ (
    .A(addr_i_5_),
    .B(_07105_),
    .C(_00498_),
    .Y(_04403_)
  );
  sg13g2_nor2_1 _14477_ (
    .A(_00297_),
    .B(_03167_),
    .Y(_04404_)
  );
  sg13g2_o21ai_1 _14478_ (
    .A1(_04403_),
    .A2(_04404_),
    .B1(addr_i_2_),
    .Y(_04405_)
  );
  sg13g2_nand2b_1 _14479_ (
    .A_N(_03039_),
    .B(_04405_),
    .Y(_04406_)
  );
  sg13g2_a22oi_1 _14480_ (
    .A1(addr_i_4_),
    .A2(_04402_),
    .B1(_04406_),
    .B2(addr_i_8_),
    .Y(_04408_)
  );
  sg13g2_a221oi_1 _14481_ (
    .A1(addr_i_8_),
    .A2(_04393_),
    .B1(_04397_),
    .B2(_04408_),
    .C1(_06652_),
    .Y(_04409_)
  );
  sg13g2_a21o_1 _14482_ (
    .A1(addr_i_3_),
    .A2(_03004_),
    .B1(_01962_),
    .X(_04410_)
  );
  sg13g2_a22oi_1 _14483_ (
    .A1(_02213_),
    .A2(_00961_),
    .B1(addr_i_2_),
    .B2(addr_i_5_),
    .Y(_04411_)
  );
  sg13g2_a22oi_1 _14484_ (
    .A1(addr_i_2_),
    .A2(_04410_),
    .B1(_04411_),
    .B2(_09271_),
    .Y(_04412_)
  );
  sg13g2_nand2_1 _14485_ (
    .A(_00484_),
    .B(_00038_),
    .Y(_04413_)
  );
  sg13g2_o21ai_1 _14486_ (
    .A1(_00700_),
    .A2(_04413_),
    .B1(_00482_),
    .Y(_04414_)
  );
  sg13g2_a22oi_1 _14487_ (
    .A1(_06619_),
    .A2(_04414_),
    .B1(_01604_),
    .B2(addr_i_4_),
    .Y(_04415_)
  );
  sg13g2_nor2_1 _14488_ (
    .A(_04412_),
    .B(_04415_),
    .Y(_04416_)
  );
  sg13g2_a22oi_1 _14489_ (
    .A1(_01437_),
    .A2(_02171_),
    .B1(_04416_),
    .B2(addr_i_8_),
    .Y(_04417_)
  );
  sg13g2_nand2_1 _14490_ (
    .A(addr_i_3_),
    .B(_01179_),
    .Y(_04419_)
  );
  sg13g2_nand2_1 _14491_ (
    .A(_00870_),
    .B(_04419_),
    .Y(_04420_)
  );
  sg13g2_nand2_1 _14492_ (
    .A(addr_i_4_),
    .B(_04420_),
    .Y(_04421_)
  );
  sg13g2_o21ai_1 _14493_ (
    .A1(_03452_),
    .A2(_03671_),
    .B1(_04421_),
    .Y(_04422_)
  );
  sg13g2_nor3_1 _14494_ (
    .A(addr_i_4_),
    .B(_08343_),
    .C(_02107_),
    .Y(_04423_)
  );
  sg13g2_a21oi_1 _14495_ (
    .A1(addr_i_5_),
    .A2(_02494_),
    .B1(_04423_),
    .Y(_04424_)
  );
  sg13g2_o21ai_1 _14496_ (
    .A1(_00053_),
    .A2(_04424_),
    .B1(addr_i_8_),
    .Y(_04425_)
  );
  sg13g2_nor2_1 _14497_ (
    .A(addr_i_5_),
    .B(_08111_),
    .Y(_04426_)
  );
  sg13g2_o21ai_1 _14498_ (
    .A1(addr_i_2_),
    .A2(_04426_),
    .B1(_05357_),
    .Y(_04427_)
  );
  sg13g2_nand2_1 _14499_ (
    .A(addr_i_6_),
    .B(_04427_),
    .Y(_04428_)
  );
  sg13g2_nor2_1 _14500_ (
    .A(_00543_),
    .B(_01432_),
    .Y(_04430_)
  );
  sg13g2_a22oi_1 _14501_ (
    .A1(_00258_),
    .A2(_09382_),
    .B1(_01846_),
    .B2(_04430_),
    .Y(_04431_)
  );
  sg13g2_a21oi_1 _14502_ (
    .A1(_04428_),
    .A2(_04431_),
    .B1(addr_i_7_),
    .Y(_04432_)
  );
  sg13g2_a22oi_1 _14503_ (
    .A1(_01892_),
    .A2(_04422_),
    .B1(_04425_),
    .B2(_04432_),
    .Y(_04433_)
  );
  sg13g2_nor3_1 _14504_ (
    .A(_00925_),
    .B(_04417_),
    .C(_04433_),
    .Y(_04434_)
  );
  sg13g2_nor4_1 _14505_ (
    .A(addr_i_11_),
    .B(_04383_),
    .C(_04409_),
    .D(_04434_),
    .Y(_04435_)
  );
  sg13g2_or3_1 _14506_ (
    .A(addr_i_12_),
    .B(_04346_),
    .C(_04435_),
    .X(_04436_)
  );
  sg13g2_o21ai_1 _14507_ (
    .A1(_04155_),
    .A2(_04258_),
    .B1(_04436_),
    .Y(data_o_20_)
  );
  sg13g2_a21oi_1 _14508_ (
    .A1(_01257_),
    .A2(_02742_),
    .B1(_02171_),
    .Y(_04437_)
  );
  sg13g2_nor3_1 _14509_ (
    .A(addr_i_4_),
    .B(_05292_),
    .C(_03984_),
    .Y(_04438_)
  );
  sg13g2_a22oi_1 _14510_ (
    .A1(addr_i_4_),
    .A2(_04437_),
    .B1(_04438_),
    .B2(addr_i_7_),
    .Y(_04440_)
  );
  sg13g2_o21ai_1 _14511_ (
    .A1(addr_i_5_),
    .A2(_01580_),
    .B1(_03577_),
    .Y(_04441_)
  );
  sg13g2_buf_1 _14512_ (
    .A(_00375_),
    .X(_04442_)
  );
  sg13g2_nand2_1 _14513_ (
    .A(_02283_),
    .B(_01199_),
    .Y(_04443_)
  );
  sg13g2_o21ai_1 _14514_ (
    .A1(_04442_),
    .A2(_00346_),
    .B1(_04443_),
    .Y(_04444_)
  );
  sg13g2_nand2_1 _14515_ (
    .A(_04441_),
    .B(_04444_),
    .Y(_04445_)
  );
  sg13g2_o21ai_1 _14516_ (
    .A1(_04440_),
    .A2(_04445_),
    .B1(_01350_),
    .Y(_04446_)
  );
  sg13g2_a21o_1 _14517_ (
    .A1(_03519_),
    .A2(_00592_),
    .B1(addr_i_4_),
    .X(_04447_)
  );
  sg13g2_o21ai_1 _14518_ (
    .A1(_00060_),
    .A2(_01697_),
    .B1(_00430_),
    .Y(_04448_)
  );
  sg13g2_o21ai_1 _14519_ (
    .A1(_08431_),
    .A2(_02578_),
    .B1(addr_i_7_),
    .Y(_04449_)
  );
  sg13g2_nand2_1 _14520_ (
    .A(_08156_),
    .B(_01033_),
    .Y(_04451_)
  );
  sg13g2_a21oi_1 _14521_ (
    .A1(_02708_),
    .A2(_04451_),
    .B1(_00146_),
    .Y(_04452_)
  );
  sg13g2_a22oi_1 _14522_ (
    .A1(addr_i_5_),
    .A2(_04448_),
    .B1(_04449_),
    .B2(_04452_),
    .Y(_04453_)
  );
  sg13g2_a21oi_1 _14523_ (
    .A1(_05834_),
    .A2(_04447_),
    .B1(_04453_),
    .Y(_04454_)
  );
  sg13g2_nor4_1 _14524_ (
    .A(_03073_),
    .B(_02536_),
    .C(_00820_),
    .D(_02179_),
    .Y(_04455_)
  );
  sg13g2_a22oi_1 _14525_ (
    .A1(_01613_),
    .A2(_04454_),
    .B1(_04455_),
    .B2(addr_i_11_),
    .Y(_04456_)
  );
  sg13g2_a221oi_1 _14526_ (
    .A1(_04442_),
    .A2(_00159_),
    .B1(_01653_),
    .B2(_01030_),
    .C1(addr_i_7_),
    .Y(_04457_)
  );
  sg13g2_o21ai_1 _14527_ (
    .A1(addr_i_4_),
    .A2(_01183_),
    .B1(_03660_),
    .Y(_04458_)
  );
  sg13g2_nand2_1 _14528_ (
    .A(addr_i_7_),
    .B(_02695_),
    .Y(_04459_)
  );
  sg13g2_a221oi_1 _14529_ (
    .A1(addr_i_3_),
    .A2(_03833_),
    .B1(_04458_),
    .B2(_00388_),
    .C1(_04459_),
    .Y(_04460_)
  );
  sg13g2_nor3_1 _14530_ (
    .A(addr_i_8_),
    .B(_04457_),
    .C(_04460_),
    .Y(_04462_)
  );
  sg13g2_nand3_1 _14531_ (
    .A(addr_i_3_),
    .B(_00186_),
    .C(_03575_),
    .Y(_04463_)
  );
  sg13g2_nor3_1 _14532_ (
    .A(addr_i_2_),
    .B(addr_i_5_),
    .C(_01319_),
    .Y(_04464_)
  );
  sg13g2_or3_1 _14533_ (
    .A(addr_i_3_),
    .B(_00946_),
    .C(_04464_),
    .X(_04465_)
  );
  sg13g2_a21oi_1 _14534_ (
    .A1(_04463_),
    .A2(_04465_),
    .B1(addr_i_4_),
    .Y(_04466_)
  );
  sg13g2_o21ai_1 _14535_ (
    .A1(_01191_),
    .A2(_09205_),
    .B1(_01060_),
    .Y(_04467_)
  );
  sg13g2_a22oi_1 _14536_ (
    .A1(_03292_),
    .A2(_04467_),
    .B1(_00026_),
    .B2(_00084_),
    .Y(_04468_)
  );
  sg13g2_nor3_1 _14537_ (
    .A(_03259_),
    .B(_04466_),
    .C(_04468_),
    .Y(_04469_)
  );
  sg13g2_o21ai_1 _14538_ (
    .A1(_04462_),
    .A2(_04469_),
    .B1(_05214_),
    .Y(_04470_)
  );
  sg13g2_nand2b_1 _14539_ (
    .A_N(_02652_),
    .B(_03248_),
    .Y(_04471_)
  );
  sg13g2_nor2_1 _14540_ (
    .A(addr_i_3_),
    .B(_00621_),
    .Y(_04473_)
  );
  sg13g2_a22oi_1 _14541_ (
    .A1(_03281_),
    .A2(_04471_),
    .B1(_04473_),
    .B2(_01528_),
    .Y(_04474_)
  );
  sg13g2_or2_1 _14542_ (
    .A(_00064_),
    .B(_02403_),
    .X(_04475_)
  );
  sg13g2_o21ai_1 _14543_ (
    .A1(addr_i_2_),
    .A2(_02761_),
    .B1(_04475_),
    .Y(_04476_)
  );
  sg13g2_a221oi_1 _14544_ (
    .A1(_08653_),
    .A2(_08188_),
    .B1(_04476_),
    .B2(addr_i_3_),
    .C1(addr_i_4_),
    .Y(_04477_)
  );
  sg13g2_nor2_1 _14545_ (
    .A(_04474_),
    .B(_04477_),
    .Y(_04478_)
  );
  sg13g2_a22oi_1 _14546_ (
    .A1(_00103_),
    .A2(_03793_),
    .B1(_04478_),
    .B2(_01043_),
    .Y(_04479_)
  );
  sg13g2_nor3_1 _14547_ (
    .A(_00381_),
    .B(_08410_),
    .C(_01747_),
    .Y(_04480_)
  );
  sg13g2_nand2_1 _14548_ (
    .A(_01972_),
    .B(_08719_),
    .Y(_04481_)
  );
  sg13g2_nor3_1 _14549_ (
    .A(_00463_),
    .B(_06143_),
    .C(_01507_),
    .Y(_04482_)
  );
  sg13g2_o21ai_1 _14550_ (
    .A1(_01652_),
    .A2(_04482_),
    .B1(addr_i_6_),
    .Y(_04484_)
  );
  sg13g2_a21oi_1 _14551_ (
    .A1(_04481_),
    .A2(_04484_),
    .B1(addr_i_4_),
    .Y(_04485_)
  );
  sg13g2_a22oi_1 _14552_ (
    .A1(_00973_),
    .A2(_04480_),
    .B1(_04485_),
    .B2(addr_i_8_),
    .Y(_04486_)
  );
  sg13g2_nor3_1 _14553_ (
    .A(addr_i_9_),
    .B(_04479_),
    .C(_04486_),
    .Y(_04487_)
  );
  sg13g2_o21ai_1 _14554_ (
    .A1(_00103_),
    .A2(_01473_),
    .B1(_01446_),
    .Y(_04488_)
  );
  sg13g2_a221oi_1 _14555_ (
    .A1(_00001_),
    .A2(_07458_),
    .B1(_00569_),
    .B2(_00959_),
    .C1(_02322_),
    .Y(_04489_)
  );
  sg13g2_nor2_1 _14556_ (
    .A(_05036_),
    .B(_00521_),
    .Y(_04490_)
  );
  sg13g2_a21oi_1 _14557_ (
    .A1(_00072_),
    .A2(_02976_),
    .B1(_04490_),
    .Y(_04491_)
  );
  sg13g2_a21oi_1 _14558_ (
    .A1(_04489_),
    .A2(_04491_),
    .B1(_02796_),
    .Y(_04492_)
  );
  sg13g2_a21oi_1 _14559_ (
    .A1(addr_i_3_),
    .A2(_04488_),
    .B1(_04492_),
    .Y(_04493_)
  );
  sg13g2_o21ai_1 _14560_ (
    .A1(addr_i_2_),
    .A2(_01033_),
    .B1(_00117_),
    .Y(_04495_)
  );
  sg13g2_nand4_1 _14561_ (
    .A(addr_i_7_),
    .B(_02920_),
    .C(_00368_),
    .D(_04495_),
    .Y(_04496_)
  );
  sg13g2_nand3_1 _14562_ (
    .A(_05811_),
    .B(_00516_),
    .C(_05612_),
    .Y(_04497_)
  );
  sg13g2_a22oi_1 _14563_ (
    .A1(_04496_),
    .A2(_04497_),
    .B1(_00565_),
    .B2(_01402_),
    .Y(_04498_)
  );
  sg13g2_nor2_1 _14564_ (
    .A(_00103_),
    .B(_00185_),
    .Y(_04499_)
  );
  sg13g2_a21oi_1 _14565_ (
    .A1(addr_i_6_),
    .A2(_01738_),
    .B1(_02479_),
    .Y(_04500_)
  );
  sg13g2_a22oi_1 _14566_ (
    .A1(_01086_),
    .A2(_01495_),
    .B1(_04500_),
    .B2(_00192_),
    .Y(_04501_)
  );
  sg13g2_nor2_1 _14567_ (
    .A(addr_i_3_),
    .B(_04501_),
    .Y(_04502_)
  );
  sg13g2_nor4_1 _14568_ (
    .A(_00629_),
    .B(_04498_),
    .C(_04499_),
    .D(_04502_),
    .Y(_04503_)
  );
  sg13g2_a22oi_1 _14569_ (
    .A1(_03259_),
    .A2(_04493_),
    .B1(_04503_),
    .B2(_00396_),
    .Y(_04504_)
  );
  sg13g2_o21ai_1 _14570_ (
    .A1(_04487_),
    .A2(_04504_),
    .B1(_00511_),
    .Y(_04507_)
  );
  sg13g2_and4_1 _14571_ (
    .A(_04446_),
    .B(_04456_),
    .C(_04470_),
    .D(_04507_),
    .X(_04508_)
  );
  sg13g2_a22oi_1 _14572_ (
    .A1(_08388_),
    .A2(_01330_),
    .B1(_01127_),
    .B2(_02327_),
    .Y(_04509_)
  );
  sg13g2_o21ai_1 _14573_ (
    .A1(_02796_),
    .A2(_04509_),
    .B1(_05611_),
    .Y(_04510_)
  );
  sg13g2_o21ai_1 _14574_ (
    .A1(_07647_),
    .A2(_08310_),
    .B1(addr_i_4_),
    .Y(_04511_)
  );
  sg13g2_o21ai_1 _14575_ (
    .A1(_01459_),
    .A2(_02774_),
    .B1(_00778_),
    .Y(_04512_)
  );
  sg13g2_nand4_1 _14576_ (
    .A(addr_i_3_),
    .B(_00138_),
    .C(_04511_),
    .D(_04512_),
    .Y(_04513_)
  );
  sg13g2_o21ai_1 _14577_ (
    .A1(addr_i_3_),
    .A2(_04510_),
    .B1(_04513_),
    .Y(_04514_)
  );
  sg13g2_a21oi_1 _14578_ (
    .A1(_04229_),
    .A2(_01740_),
    .B1(addr_i_6_),
    .Y(_04515_)
  );
  sg13g2_nor2_1 _14579_ (
    .A(_02700_),
    .B(_04515_),
    .Y(_04516_)
  );
  sg13g2_o21ai_1 _14580_ (
    .A1(_00783_),
    .A2(_02171_),
    .B1(_00268_),
    .Y(_04518_)
  );
  sg13g2_o21ai_1 _14581_ (
    .A1(_01015_),
    .A2(_05932_),
    .B1(addr_i_3_),
    .Y(_04519_)
  );
  sg13g2_nand2_1 _14582_ (
    .A(_04518_),
    .B(_04519_),
    .Y(_04520_)
  );
  sg13g2_nor2_1 _14583_ (
    .A(_00799_),
    .B(_02055_),
    .Y(_04521_)
  );
  sg13g2_a22oi_1 _14584_ (
    .A1(addr_i_4_),
    .A2(_02166_),
    .B1(_01500_),
    .B2(addr_i_3_),
    .Y(_04522_)
  );
  sg13g2_a22oi_1 _14585_ (
    .A1(_02956_),
    .A2(_04521_),
    .B1(_04522_),
    .B2(addr_i_7_),
    .Y(_04523_)
  );
  sg13g2_a22oi_1 _14586_ (
    .A1(addr_i_7_),
    .A2(_04520_),
    .B1(_04523_),
    .B2(addr_i_9_),
    .Y(_04524_)
  );
  sg13g2_a22oi_1 _14587_ (
    .A1(_04514_),
    .A2(_04516_),
    .B1(_04524_),
    .B2(addr_i_8_),
    .Y(_04525_)
  );
  sg13g2_o21ai_1 _14588_ (
    .A1(_01015_),
    .A2(_00192_),
    .B1(addr_i_3_),
    .Y(_04526_)
  );
  sg13g2_nand2b_1 _14589_ (
    .A_N(_06519_),
    .B(_04526_),
    .Y(_04527_)
  );
  sg13g2_nand2_1 _14590_ (
    .A(_03964_),
    .B(_01420_),
    .Y(_04529_)
  );
  sg13g2_a21oi_1 _14591_ (
    .A1(_01594_),
    .A2(_04529_),
    .B1(addr_i_3_),
    .Y(_04530_)
  );
  sg13g2_a21oi_1 _14592_ (
    .A1(_00926_),
    .A2(_01661_),
    .B1(addr_i_6_),
    .Y(_04531_)
  );
  sg13g2_a22oi_1 _14593_ (
    .A1(addr_i_7_),
    .A2(_04527_),
    .B1(_04530_),
    .B2(_04531_),
    .Y(_04532_)
  );
  sg13g2_o21ai_1 _14594_ (
    .A1(_01439_),
    .A2(_02848_),
    .B1(addr_i_2_),
    .Y(_04533_)
  );
  sg13g2_nand3_1 _14595_ (
    .A(addr_i_3_),
    .B(addr_i_7_),
    .C(_00566_),
    .Y(_04534_)
  );
  sg13g2_nand3_1 _14596_ (
    .A(addr_i_4_),
    .B(_04533_),
    .C(_04534_),
    .Y(_04535_)
  );
  sg13g2_nand2b_1 _14597_ (
    .A_N(_01808_),
    .B(_01946_),
    .Y(_04536_)
  );
  sg13g2_nand3_1 _14598_ (
    .A(addr_i_3_),
    .B(_00056_),
    .C(_00453_),
    .Y(_04537_)
  );
  sg13g2_nor2_1 _14599_ (
    .A(_00624_),
    .B(_00676_),
    .Y(_04538_)
  );
  sg13g2_nand2_1 _14600_ (
    .A(_08000_),
    .B(_04538_),
    .Y(_04540_)
  );
  sg13g2_nand3_1 _14601_ (
    .A(_00910_),
    .B(_01155_),
    .C(_04540_),
    .Y(_04541_)
  );
  sg13g2_nand3_1 _14602_ (
    .A(addr_i_9_),
    .B(addr_i_8_),
    .C(_01441_),
    .Y(_04542_)
  );
  sg13g2_a221oi_1 _14603_ (
    .A1(_04535_),
    .A2(_04536_),
    .B1(_04537_),
    .B2(_04541_),
    .C1(_04542_),
    .Y(_04543_)
  );
  sg13g2_nor2_1 _14604_ (
    .A(addr_i_10_),
    .B(_04543_),
    .Y(_04544_)
  );
  sg13g2_o21ai_1 _14605_ (
    .A1(_01612_),
    .A2(_04532_),
    .B1(_04544_),
    .Y(_04545_)
  );
  sg13g2_o21ai_1 _14606_ (
    .A1(_00298_),
    .A2(_00597_),
    .B1(_00565_),
    .Y(_04546_)
  );
  sg13g2_a21oi_1 _14607_ (
    .A1(_00785_),
    .A2(_04252_),
    .B1(_00046_),
    .Y(_04547_)
  );
  sg13g2_o21ai_1 _14608_ (
    .A1(_02203_),
    .A2(_04547_),
    .B1(_02344_),
    .Y(_04548_)
  );
  sg13g2_a21oi_1 _14609_ (
    .A1(_00566_),
    .A2(_00470_),
    .B1(_00648_),
    .Y(_04549_)
  );
  sg13g2_o21ai_1 _14610_ (
    .A1(_00205_),
    .A2(_04549_),
    .B1(addr_i_2_),
    .Y(_04551_)
  );
  sg13g2_nand4_1 _14611_ (
    .A(addr_i_7_),
    .B(_04546_),
    .C(_04548_),
    .D(_04551_),
    .Y(_04552_)
  );
  sg13g2_nor2_1 _14612_ (
    .A(_09510_),
    .B(_07911_),
    .Y(_04553_)
  );
  sg13g2_a22oi_1 _14613_ (
    .A1(_00990_),
    .A2(_07911_),
    .B1(_04553_),
    .B2(addr_i_4_),
    .Y(_04554_)
  );
  sg13g2_a21oi_1 _14614_ (
    .A1(_00482_),
    .A2(_09415_),
    .B1(addr_i_3_),
    .Y(_04555_)
  );
  sg13g2_nor3_1 _14615_ (
    .A(_01131_),
    .B(_03742_),
    .C(_04555_),
    .Y(_04556_)
  );
  sg13g2_o21ai_1 _14616_ (
    .A1(_04554_),
    .A2(_04556_),
    .B1(_01475_),
    .Y(_04557_)
  );
  sg13g2_nand3_1 _14617_ (
    .A(_00423_),
    .B(_04552_),
    .C(_04557_),
    .Y(_04558_)
  );
  sg13g2_nand2_1 _14618_ (
    .A(_00967_),
    .B(_04213_),
    .Y(_04559_)
  );
  sg13g2_nor2_1 _14619_ (
    .A(_02063_),
    .B(_00132_),
    .Y(_04560_)
  );
  sg13g2_a22oi_1 _14620_ (
    .A1(_00183_),
    .A2(_01367_),
    .B1(_00087_),
    .B2(addr_i_5_),
    .Y(_04562_)
  );
  sg13g2_a22oi_1 _14621_ (
    .A1(_04559_),
    .A2(_04560_),
    .B1(_04562_),
    .B2(_01935_),
    .Y(_04563_)
  );
  sg13g2_mux2_1 _14622_ (
    .A0(_01622_),
    .A1(_03631_),
    .S(addr_i_4_),
    .X(_04564_)
  );
  sg13g2_nor2_1 _14623_ (
    .A(_02472_),
    .B(_01949_),
    .Y(_04565_)
  );
  sg13g2_a21oi_1 _14624_ (
    .A1(addr_i_2_),
    .A2(_04564_),
    .B1(_04565_),
    .Y(_04566_)
  );
  sg13g2_nand2_1 _14625_ (
    .A(_00298_),
    .B(_09499_),
    .Y(_04567_)
  );
  sg13g2_o21ai_1 _14626_ (
    .A1(addr_i_3_),
    .A2(_04566_),
    .B1(_04567_),
    .Y(_04568_)
  );
  sg13g2_o21ai_1 _14627_ (
    .A1(_04563_),
    .A2(_04568_),
    .B1(_02604_),
    .Y(_04569_)
  );
  sg13g2_o21ai_1 _14628_ (
    .A1(_00569_),
    .A2(_01845_),
    .B1(_00168_),
    .Y(_04570_)
  );
  sg13g2_o21ai_1 _14629_ (
    .A1(_02479_),
    .A2(_02107_),
    .B1(_02656_),
    .Y(_04571_)
  );
  sg13g2_a22oi_1 _14630_ (
    .A1(_02470_),
    .A2(_00543_),
    .B1(_00844_),
    .B2(_02569_),
    .Y(_04573_)
  );
  sg13g2_a22oi_1 _14631_ (
    .A1(_05247_),
    .A2(_04571_),
    .B1(_04573_),
    .B2(_07282_),
    .Y(_04574_)
  );
  sg13g2_a21oi_1 _14632_ (
    .A1(_02250_),
    .A2(_03845_),
    .B1(addr_i_3_),
    .Y(_04575_)
  );
  sg13g2_o21ai_1 _14633_ (
    .A1(_02801_),
    .A2(_04575_),
    .B1(_00262_),
    .Y(_04576_)
  );
  sg13g2_nand3_1 _14634_ (
    .A(_04570_),
    .B(_04574_),
    .C(_04576_),
    .Y(_04577_)
  );
  sg13g2_a21oi_1 _14635_ (
    .A1(_00736_),
    .A2(_05457_),
    .B1(_05711_),
    .Y(_04578_)
  );
  sg13g2_nand2_1 _14636_ (
    .A(addr_i_2_),
    .B(_00380_),
    .Y(_04579_)
  );
  sg13g2_a21oi_1 _14637_ (
    .A1(_00831_),
    .A2(_04579_),
    .B1(addr_i_3_),
    .Y(_04580_)
  );
  sg13g2_o21ai_1 _14638_ (
    .A1(_04578_),
    .A2(_04580_),
    .B1(_01878_),
    .Y(_04581_)
  );
  sg13g2_o21ai_1 _14639_ (
    .A1(_06298_),
    .A2(_01107_),
    .B1(addr_i_3_),
    .Y(_04582_)
  );
  sg13g2_a22oi_1 _14640_ (
    .A1(_06607_),
    .A2(_00727_),
    .B1(_06563_),
    .B2(_05811_),
    .Y(_04584_)
  );
  sg13g2_nand3_1 _14641_ (
    .A(addr_i_3_),
    .B(_00581_),
    .C(_01636_),
    .Y(_04585_)
  );
  sg13g2_a21oi_1 _14642_ (
    .A1(_02864_),
    .A2(_04585_),
    .B1(_02294_),
    .Y(_04586_)
  );
  sg13g2_a22oi_1 _14643_ (
    .A1(_04582_),
    .A2(_04584_),
    .B1(_04586_),
    .B2(addr_i_8_),
    .Y(_04587_)
  );
  sg13g2_a21oi_1 _14644_ (
    .A1(_04581_),
    .A2(_04587_),
    .B1(_09315_),
    .Y(_04588_)
  );
  sg13g2_nand2_1 _14645_ (
    .A(_04577_),
    .B(_04588_),
    .Y(_04589_)
  );
  sg13g2_nand4_1 _14646_ (
    .A(addr_i_10_),
    .B(_04558_),
    .C(_04569_),
    .D(_04589_),
    .Y(_04590_)
  );
  sg13g2_o21ai_1 _14647_ (
    .A1(_04525_),
    .A2(_04545_),
    .B1(_04590_),
    .Y(_04591_)
  );
  sg13g2_a21o_1 _14648_ (
    .A1(addr_i_11_),
    .A2(_04591_),
    .B1(addr_i_12_),
    .X(_04592_)
  );
  sg13g2_o21ai_1 _14649_ (
    .A1(_01380_),
    .A2(_03577_),
    .B1(addr_i_3_),
    .Y(_04593_)
  );
  sg13g2_a21oi_1 _14650_ (
    .A1(_00567_),
    .A2(_00671_),
    .B1(addr_i_3_),
    .Y(_04595_)
  );
  sg13g2_nor4_1 _14651_ (
    .A(_04068_),
    .B(_02265_),
    .C(_03565_),
    .D(_04595_),
    .Y(_04596_)
  );
  sg13g2_o21ai_1 _14652_ (
    .A1(_02479_),
    .A2(_08774_),
    .B1(_02930_),
    .Y(_04597_)
  );
  sg13g2_a22oi_1 _14653_ (
    .A1(addr_i_3_),
    .A2(_04597_),
    .B1(_02374_),
    .B2(addr_i_7_),
    .Y(_04598_)
  );
  sg13g2_a22oi_1 _14654_ (
    .A1(_04593_),
    .A2(_04596_),
    .B1(_04598_),
    .B2(_00214_),
    .Y(_04599_)
  );
  sg13g2_o21ai_1 _14655_ (
    .A1(_08166_),
    .A2(_00494_),
    .B1(addr_i_2_),
    .Y(_04600_)
  );
  sg13g2_o21ai_1 _14656_ (
    .A1(addr_i_3_),
    .A2(_09215_),
    .B1(_04600_),
    .Y(_04601_)
  );
  sg13g2_a221oi_1 _14657_ (
    .A1(_01019_),
    .A2(_02567_),
    .B1(_04601_),
    .B2(addr_i_6_),
    .C1(addr_i_7_),
    .Y(_04602_)
  );
  sg13g2_nor3_1 _14658_ (
    .A(_01611_),
    .B(_03631_),
    .C(_04602_),
    .Y(_04603_)
  );
  sg13g2_nand2_1 _14659_ (
    .A(_01310_),
    .B(_00972_),
    .Y(_04604_)
  );
  sg13g2_o21ai_1 _14660_ (
    .A1(_01666_),
    .A2(_00666_),
    .B1(_04604_),
    .Y(_04606_)
  );
  sg13g2_nor2_1 _14661_ (
    .A(_02700_),
    .B(_04606_),
    .Y(_04607_)
  );
  sg13g2_or3_1 _14662_ (
    .A(_04599_),
    .B(_04603_),
    .C(_04607_),
    .X(_04608_)
  );
  sg13g2_a21oi_1 _14663_ (
    .A1(_04439_),
    .A2(_07558_),
    .B1(_01645_),
    .Y(_04609_)
  );
  sg13g2_o21ai_1 _14664_ (
    .A1(_02040_),
    .A2(_04609_),
    .B1(addr_i_11_),
    .Y(_04610_)
  );
  sg13g2_a21o_1 _14665_ (
    .A1(_01774_),
    .A2(_04608_),
    .B1(_04610_),
    .X(_04611_)
  );
  sg13g2_a21oi_1 _14666_ (
    .A1(_02107_),
    .A2(_00578_),
    .B1(_00839_),
    .Y(_04612_)
  );
  sg13g2_nor2_1 _14667_ (
    .A(_03765_),
    .B(_00577_),
    .Y(_04613_)
  );
  sg13g2_o21ai_1 _14668_ (
    .A1(_02015_),
    .A2(_04613_),
    .B1(_01308_),
    .Y(_04614_)
  );
  sg13g2_o21ai_1 _14669_ (
    .A1(addr_i_5_),
    .A2(_04612_),
    .B1(_04614_),
    .Y(_04615_)
  );
  sg13g2_nor2_1 _14670_ (
    .A(_00483_),
    .B(_00557_),
    .Y(_04618_)
  );
  sg13g2_nand2_1 _14671_ (
    .A(_00704_),
    .B(_04618_),
    .Y(_04619_)
  );
  sg13g2_o21ai_1 _14672_ (
    .A1(_08896_),
    .A2(_00011_),
    .B1(_00354_),
    .Y(_04620_)
  );
  sg13g2_nand3_1 _14673_ (
    .A(_01674_),
    .B(_01257_),
    .C(_04620_),
    .Y(_04621_)
  );
  sg13g2_a21oi_1 _14674_ (
    .A1(_02815_),
    .A2(_08951_),
    .B1(_00261_),
    .Y(_04622_)
  );
  sg13g2_a22oi_1 _14675_ (
    .A1(_04619_),
    .A2(_04621_),
    .B1(_04622_),
    .B2(_03227_),
    .Y(_04623_)
  );
  sg13g2_o21ai_1 _14676_ (
    .A1(_02424_),
    .A2(_09348_),
    .B1(addr_i_3_),
    .Y(_04624_)
  );
  sg13g2_a21oi_1 _14677_ (
    .A1(addr_i_4_),
    .A2(_03458_),
    .B1(_01274_),
    .Y(_04625_)
  );
  sg13g2_nand2_1 _14678_ (
    .A(_04624_),
    .B(_04625_),
    .Y(_04626_)
  );
  sg13g2_a21oi_1 _14679_ (
    .A1(_01813_),
    .A2(_02507_),
    .B1(addr_i_3_),
    .Y(_04627_)
  );
  sg13g2_o21ai_1 _14680_ (
    .A1(_04626_),
    .A2(_04627_),
    .B1(addr_i_9_),
    .Y(_04629_)
  );
  sg13g2_a22oi_1 _14681_ (
    .A1(_00610_),
    .A2(_04615_),
    .B1(_04623_),
    .B2(_04629_),
    .Y(_04630_)
  );
  sg13g2_nor3_1 _14682_ (
    .A(addr_i_3_),
    .B(addr_i_5_),
    .C(_08763_),
    .Y(_04631_)
  );
  sg13g2_nand2_1 _14683_ (
    .A(addr_i_3_),
    .B(_07636_),
    .Y(_04632_)
  );
  sg13g2_a21oi_1 _14684_ (
    .A1(_01077_),
    .A2(_04632_),
    .B1(_00293_),
    .Y(_04633_)
  );
  sg13g2_o21ai_1 _14685_ (
    .A1(_04631_),
    .A2(_04633_),
    .B1(addr_i_4_),
    .Y(_04634_)
  );
  sg13g2_o21ai_1 _14686_ (
    .A1(_09459_),
    .A2(_00945_),
    .B1(_01302_),
    .Y(_04635_)
  );
  sg13g2_a21o_1 _14687_ (
    .A1(_04634_),
    .A2(_04635_),
    .B1(_07614_),
    .X(_04636_)
  );
  sg13g2_a21oi_1 _14688_ (
    .A1(_04893_),
    .A2(_01524_),
    .B1(_00956_),
    .Y(_04637_)
  );
  sg13g2_a21oi_1 _14689_ (
    .A1(_02369_),
    .A2(_01493_),
    .B1(_04637_),
    .Y(_04638_)
  );
  sg13g2_nand2_1 _14690_ (
    .A(_09501_),
    .B(_05424_),
    .Y(_04640_)
  );
  sg13g2_o21ai_1 _14691_ (
    .A1(_00521_),
    .A2(_00299_),
    .B1(_04640_),
    .Y(_04641_)
  );
  sg13g2_nor2_1 _14692_ (
    .A(_00498_),
    .B(_01152_),
    .Y(_04642_)
  );
  sg13g2_a21oi_1 _14693_ (
    .A1(addr_i_2_),
    .A2(_04641_),
    .B1(_04642_),
    .Y(_04643_)
  );
  sg13g2_o21ai_1 _14694_ (
    .A1(addr_i_2_),
    .A2(_04638_),
    .B1(_04643_),
    .Y(_04644_)
  );
  sg13g2_a21oi_1 _14695_ (
    .A1(_04760_),
    .A2(_02822_),
    .B1(addr_i_3_),
    .Y(_04645_)
  );
  sg13g2_a21oi_1 _14696_ (
    .A1(_00370_),
    .A2(_00894_),
    .B1(addr_i_7_),
    .Y(_04646_)
  );
  sg13g2_a22oi_1 _14697_ (
    .A1(_01202_),
    .A2(_08553_),
    .B1(_04646_),
    .B2(addr_i_8_),
    .Y(_04647_)
  );
  sg13g2_nor2b_1 _14698_ (
    .A(_04645_),
    .B_N(_04647_),
    .Y(_04648_)
  );
  sg13g2_a21oi_1 _14699_ (
    .A1(_00032_),
    .A2(_00719_),
    .B1(addr_i_2_),
    .Y(_04649_)
  );
  sg13g2_a21oi_1 _14700_ (
    .A1(_00927_),
    .A2(_00482_),
    .B1(_01970_),
    .Y(_04651_)
  );
  sg13g2_o21ai_1 _14701_ (
    .A1(_04649_),
    .A2(_04651_),
    .B1(addr_i_4_),
    .Y(_04652_)
  );
  sg13g2_a221oi_1 _14702_ (
    .A1(addr_i_8_),
    .A2(_04644_),
    .B1(_04648_),
    .B2(_04652_),
    .C1(addr_i_9_),
    .Y(_04653_)
  );
  sg13g2_a22oi_1 _14703_ (
    .A1(_04630_),
    .A2(_04636_),
    .B1(_04653_),
    .B2(addr_i_10_),
    .Y(_04654_)
  );
  sg13g2_nand2_1 _14704_ (
    .A(_00566_),
    .B(_00413_),
    .Y(_04655_)
  );
  sg13g2_a22oi_1 _14705_ (
    .A1(addr_i_3_),
    .A2(_04655_),
    .B1(_03858_),
    .B2(_07425_),
    .Y(_04656_)
  );
  sg13g2_nor2_1 _14706_ (
    .A(_02803_),
    .B(_04656_),
    .Y(_04657_)
  );
  sg13g2_nor2_1 _14707_ (
    .A(_01292_),
    .B(_07647_),
    .Y(_04658_)
  );
  sg13g2_a22oi_1 _14708_ (
    .A1(addr_i_3_),
    .A2(_04658_),
    .B1(_03300_),
    .B2(addr_i_4_),
    .Y(_04659_)
  );
  sg13g2_o21ai_1 _14709_ (
    .A1(_04657_),
    .A2(_04659_),
    .B1(_00708_),
    .Y(_04660_)
  );
  sg13g2_nand2_1 _14710_ (
    .A(_01113_),
    .B(_00664_),
    .Y(_04662_)
  );
  sg13g2_o21ai_1 _14711_ (
    .A1(_00442_),
    .A2(_03720_),
    .B1(addr_i_2_),
    .Y(_04663_)
  );
  sg13g2_nand2_1 _14712_ (
    .A(_06054_),
    .B(_00904_),
    .Y(_04664_)
  );
  sg13g2_o21ai_1 _14713_ (
    .A1(_00557_),
    .A2(_01112_),
    .B1(_07458_),
    .Y(_04665_)
  );
  sg13g2_nand4_1 _14714_ (
    .A(_04662_),
    .B(_04663_),
    .C(_04664_),
    .D(_04665_),
    .Y(_04666_)
  );
  sg13g2_a22oi_1 _14715_ (
    .A1(addr_i_3_),
    .A2(_02785_),
    .B1(_00839_),
    .B2(_04539_),
    .Y(_04667_)
  );
  sg13g2_o21ai_1 _14716_ (
    .A1(_06054_),
    .A2(_00177_),
    .B1(_00091_),
    .Y(_04668_)
  );
  sg13g2_o21ai_1 _14717_ (
    .A1(addr_i_5_),
    .A2(_04667_),
    .B1(_04668_),
    .Y(_04669_)
  );
  sg13g2_nand2_1 _14718_ (
    .A(_01872_),
    .B(_01453_),
    .Y(_04670_)
  );
  sg13g2_nand2_1 _14719_ (
    .A(_05711_),
    .B(_02626_),
    .Y(_04671_)
  );
  sg13g2_a21oi_1 _14720_ (
    .A1(_04419_),
    .A2(_04671_),
    .B1(addr_i_4_),
    .Y(_04673_)
  );
  sg13g2_o21ai_1 _14721_ (
    .A1(_06398_),
    .A2(_01472_),
    .B1(_02387_),
    .Y(_04674_)
  );
  sg13g2_nand3_1 _14722_ (
    .A(_00429_),
    .B(_02052_),
    .C(_04674_),
    .Y(_04675_)
  );
  sg13g2_a22oi_1 _14723_ (
    .A1(addr_i_6_),
    .A2(_04670_),
    .B1(_04673_),
    .B2(_04675_),
    .Y(_04676_)
  );
  sg13g2_a221oi_1 _14724_ (
    .A1(_00276_),
    .A2(_04666_),
    .B1(_04669_),
    .B2(_01666_),
    .C1(_04676_),
    .Y(_04677_)
  );
  sg13g2_a21oi_1 _14725_ (
    .A1(_04660_),
    .A2(_04677_),
    .B1(_06652_),
    .Y(_04678_)
  );
  sg13g2_nor2_1 _14726_ (
    .A(_01729_),
    .B(_00543_),
    .Y(_04679_)
  );
  sg13g2_o21ai_1 _14727_ (
    .A1(_06497_),
    .A2(_02935_),
    .B1(addr_i_4_),
    .Y(_04680_)
  );
  sg13g2_nor2_1 _14728_ (
    .A(_00413_),
    .B(_00521_),
    .Y(_04681_)
  );
  sg13g2_a21oi_1 _14729_ (
    .A1(_01077_),
    .A2(_03167_),
    .B1(_00700_),
    .Y(_04682_)
  );
  sg13g2_o21ai_1 _14730_ (
    .A1(_04681_),
    .A2(_04682_),
    .B1(addr_i_5_),
    .Y(_04684_)
  );
  sg13g2_nand3b_1 _14731_ (
    .A_N(_04679_),
    .B(_04680_),
    .C(_04684_),
    .Y(_04685_)
  );
  sg13g2_nand2_1 _14732_ (
    .A(_06630_),
    .B(_04685_),
    .Y(_04686_)
  );
  sg13g2_a22oi_1 _14733_ (
    .A1(addr_i_3_),
    .A2(_02560_),
    .B1(_01041_),
    .B2(_07889_),
    .Y(_04687_)
  );
  sg13g2_nor3_1 _14734_ (
    .A(_00548_),
    .B(_00315_),
    .C(_00844_),
    .Y(_04688_)
  );
  sg13g2_a22oi_1 _14735_ (
    .A1(_00169_),
    .A2(_04687_),
    .B1(_04688_),
    .B2(addr_i_8_),
    .Y(_04689_)
  );
  sg13g2_a21oi_1 _14736_ (
    .A1(_00582_),
    .A2(_01203_),
    .B1(addr_i_3_),
    .Y(_04690_)
  );
  sg13g2_a21o_1 _14737_ (
    .A1(_00542_),
    .A2(_06983_),
    .B1(_04690_),
    .X(_04691_)
  );
  sg13g2_o21ai_1 _14738_ (
    .A1(_04539_),
    .A2(_01954_),
    .B1(addr_i_7_),
    .Y(_04692_)
  );
  sg13g2_nor2_1 _14739_ (
    .A(_02196_),
    .B(_00384_),
    .Y(_04693_)
  );
  sg13g2_o21ai_1 _14740_ (
    .A1(_08575_),
    .A2(_04693_),
    .B1(addr_i_5_),
    .Y(_04695_)
  );
  sg13g2_a21oi_1 _14741_ (
    .A1(_00260_),
    .A2(_06972_),
    .B1(addr_i_4_),
    .Y(_04696_)
  );
  sg13g2_o21ai_1 _14742_ (
    .A1(_00977_),
    .A2(_04696_),
    .B1(addr_i_3_),
    .Y(_04697_)
  );
  sg13g2_and4_1 _14743_ (
    .A(_02027_),
    .B(_04692_),
    .C(_04695_),
    .D(_04697_),
    .X(_04698_)
  );
  sg13g2_o21ai_1 _14744_ (
    .A1(_08056_),
    .A2(_06950_),
    .B1(_00159_),
    .Y(_04699_)
  );
  sg13g2_nand3_1 _14745_ (
    .A(_00168_),
    .B(_00607_),
    .C(_02536_),
    .Y(_04700_)
  );
  sg13g2_nand3_1 _14746_ (
    .A(addr_i_8_),
    .B(_04699_),
    .C(_04700_),
    .Y(_04701_)
  );
  sg13g2_a22oi_1 _14747_ (
    .A1(addr_i_6_),
    .A2(_04691_),
    .B1(_04698_),
    .B2(_04701_),
    .Y(_04702_)
  );
  sg13g2_a22oi_1 _14748_ (
    .A1(_04686_),
    .A2(_04689_),
    .B1(_04702_),
    .B2(_02221_),
    .Y(_04703_)
  );
  sg13g2_or4_1 _14749_ (
    .A(addr_i_11_),
    .B(_04654_),
    .C(_04678_),
    .D(_04703_),
    .X(_04704_)
  );
  sg13g2_nand3_1 _14750_ (
    .A(addr_i_12_),
    .B(_04611_),
    .C(_04704_),
    .Y(_04706_)
  );
  sg13g2_o21ai_1 _14751_ (
    .A1(_04508_),
    .A2(_04592_),
    .B1(_04706_),
    .Y(data_o_21_)
  );
  sg13g2_nor3_1 _14752_ (
    .A(addr_i_6_),
    .B(_07270_),
    .C(_00279_),
    .Y(_04707_)
  );
  sg13g2_nor2_1 _14753_ (
    .A(_00822_),
    .B(_03761_),
    .Y(_04708_)
  );
  sg13g2_nor2_1 _14754_ (
    .A(_04707_),
    .B(_04708_),
    .Y(_04709_)
  );
  sg13g2_a21oi_1 _14755_ (
    .A1(_00749_),
    .A2(_02832_),
    .B1(_00967_),
    .Y(_04710_)
  );
  sg13g2_nor2_1 _14756_ (
    .A(_02361_),
    .B(_04710_),
    .Y(_04711_)
  );
  sg13g2_o21ai_1 _14757_ (
    .A1(addr_i_4_),
    .A2(_04709_),
    .B1(_04711_),
    .Y(_04712_)
  );
  sg13g2_nand2_1 _14758_ (
    .A(_02832_),
    .B(_00719_),
    .Y(_04713_)
  );
  sg13g2_a21o_1 _14759_ (
    .A1(addr_i_4_),
    .A2(_04713_),
    .B1(_03455_),
    .X(_04714_)
  );
  sg13g2_nor2_1 _14760_ (
    .A(_03033_),
    .B(_01227_),
    .Y(_04716_)
  );
  sg13g2_o21ai_1 _14761_ (
    .A1(_04396_),
    .A2(_04716_),
    .B1(addr_i_8_),
    .Y(_04717_)
  );
  sg13g2_a221oi_1 _14762_ (
    .A1(addr_i_7_),
    .A2(_04712_),
    .B1(_04714_),
    .B2(_09487_),
    .C1(_04717_),
    .Y(_04718_)
  );
  sg13g2_o21ai_1 _14763_ (
    .A1(_07625_),
    .A2(_07050_),
    .B1(_00677_),
    .Y(_04719_)
  );
  sg13g2_mux2_1 _14764_ (
    .A0(_04284_),
    .A1(_09485_),
    .S(addr_i_4_),
    .X(_04720_)
  );
  sg13g2_nor2_1 _14765_ (
    .A(_02744_),
    .B(_00056_),
    .Y(_04721_)
  );
  sg13g2_a21oi_1 _14766_ (
    .A1(_01480_),
    .A2(_04720_),
    .B1(_04721_),
    .Y(_04722_)
  );
  sg13g2_o21ai_1 _14767_ (
    .A1(_01155_),
    .A2(_00972_),
    .B1(_01692_),
    .Y(_04723_)
  );
  sg13g2_nor2_1 _14768_ (
    .A(_07911_),
    .B(_00660_),
    .Y(_04724_)
  );
  sg13g2_a22oi_1 _14769_ (
    .A1(_01336_),
    .A2(_04723_),
    .B1(_04724_),
    .B2(addr_i_8_),
    .Y(_04725_)
  );
  sg13g2_o21ai_1 _14770_ (
    .A1(addr_i_2_),
    .A2(_04722_),
    .B1(_04725_),
    .Y(_04728_)
  );
  sg13g2_a21oi_1 _14771_ (
    .A1(addr_i_3_),
    .A2(_04719_),
    .B1(_04728_),
    .Y(_04729_)
  );
  sg13g2_nor3_1 _14772_ (
    .A(_00109_),
    .B(_04718_),
    .C(_04729_),
    .Y(_04730_)
  );
  sg13g2_nand2_1 _14773_ (
    .A(_04672_),
    .B(_00688_),
    .Y(_04731_)
  );
  sg13g2_o21ai_1 _14774_ (
    .A1(_02501_),
    .A2(_00401_),
    .B1(_04731_),
    .Y(_04732_)
  );
  sg13g2_a22oi_1 _14775_ (
    .A1(addr_i_3_),
    .A2(_04732_),
    .B1(_00844_),
    .B2(_00507_),
    .Y(_04733_)
  );
  sg13g2_a21oi_1 _14776_ (
    .A1(_01047_),
    .A2(_01782_),
    .B1(_00717_),
    .Y(_04734_)
  );
  sg13g2_nand2_1 _14777_ (
    .A(addr_i_2_),
    .B(_04734_),
    .Y(_04735_)
  );
  sg13g2_o21ai_1 _14778_ (
    .A1(addr_i_2_),
    .A2(_04733_),
    .B1(_04735_),
    .Y(_04736_)
  );
  sg13g2_o21ai_1 _14779_ (
    .A1(_02639_),
    .A2(_00132_),
    .B1(addr_i_2_),
    .Y(_04737_)
  );
  sg13g2_o21ai_1 _14780_ (
    .A1(_00096_),
    .A2(_01567_),
    .B1(addr_i_3_),
    .Y(_04739_)
  );
  sg13g2_o21ai_1 _14781_ (
    .A1(addr_i_3_),
    .A2(_04737_),
    .B1(_04739_),
    .Y(_04740_)
  );
  sg13g2_nand2_1 _14782_ (
    .A(_00383_),
    .B(_03676_),
    .Y(_04741_)
  );
  sg13g2_o21ai_1 _14783_ (
    .A1(_01232_),
    .A2(_02632_),
    .B1(addr_i_3_),
    .Y(_04742_)
  );
  sg13g2_a21oi_1 _14784_ (
    .A1(_04741_),
    .A2(_04742_),
    .B1(addr_i_2_),
    .Y(_04743_)
  );
  sg13g2_a21o_1 _14785_ (
    .A1(addr_i_5_),
    .A2(_04740_),
    .B1(_04743_),
    .X(_04744_)
  );
  sg13g2_nand3_1 _14786_ (
    .A(_00497_),
    .B(_01462_),
    .C(_01463_),
    .Y(_04745_)
  );
  sg13g2_a21oi_1 _14787_ (
    .A1(_02820_),
    .A2(_04745_),
    .B1(_01663_),
    .Y(_04746_)
  );
  sg13g2_nor2_1 _14788_ (
    .A(_09493_),
    .B(_01022_),
    .Y(_04747_)
  );
  sg13g2_nand2_1 _14789_ (
    .A(addr_i_2_),
    .B(_07934_),
    .Y(_04748_)
  );
  sg13g2_a22oi_1 _14790_ (
    .A1(addr_i_3_),
    .A2(_04747_),
    .B1(_04748_),
    .B2(_03364_),
    .Y(_04750_)
  );
  sg13g2_nor3_1 _14791_ (
    .A(_09105_),
    .B(_00712_),
    .C(_03132_),
    .Y(_04751_)
  );
  sg13g2_or3_1 _14792_ (
    .A(addr_i_9_),
    .B(_04750_),
    .C(_04751_),
    .X(_04752_)
  );
  sg13g2_a22oi_1 _14793_ (
    .A1(_00114_),
    .A2(_04744_),
    .B1(_04746_),
    .B2(_04752_),
    .Y(_04753_)
  );
  sg13g2_nand2_1 _14794_ (
    .A(addr_i_3_),
    .B(_09371_),
    .Y(_04754_)
  );
  sg13g2_o21ai_1 _14795_ (
    .A1(addr_i_6_),
    .A2(_00818_),
    .B1(_02742_),
    .Y(_04755_)
  );
  sg13g2_nand2_1 _14796_ (
    .A(_01633_),
    .B(_04755_),
    .Y(_04756_)
  );
  sg13g2_a21oi_1 _14797_ (
    .A1(_02815_),
    .A2(_00687_),
    .B1(addr_i_3_),
    .Y(_04757_)
  );
  sg13g2_a22oi_1 _14798_ (
    .A1(_00084_),
    .A2(_04754_),
    .B1(_04756_),
    .B2(_04757_),
    .Y(_04758_)
  );
  sg13g2_or3_1 _14799_ (
    .A(_08575_),
    .B(_01025_),
    .C(_01016_),
    .X(_04759_)
  );
  sg13g2_a21oi_1 _14800_ (
    .A1(_02297_),
    .A2(_02930_),
    .B1(_08266_),
    .Y(_04761_)
  );
  sg13g2_a22oi_1 _14801_ (
    .A1(addr_i_5_),
    .A2(_04759_),
    .B1(_04761_),
    .B2(_01031_),
    .Y(_04762_)
  );
  sg13g2_nor2_1 _14802_ (
    .A(_03062_),
    .B(_04762_),
    .Y(_04763_)
  );
  sg13g2_nand2_1 _14803_ (
    .A(_00371_),
    .B(_01367_),
    .Y(_04764_)
  );
  sg13g2_o21ai_1 _14804_ (
    .A1(_02108_),
    .A2(_00303_),
    .B1(addr_i_3_),
    .Y(_04765_)
  );
  sg13g2_a21oi_1 _14805_ (
    .A1(_00567_),
    .A2(_04765_),
    .B1(addr_i_2_),
    .Y(_04766_)
  );
  sg13g2_nand2_1 _14806_ (
    .A(addr_i_7_),
    .B(_02810_),
    .Y(_04767_)
  );
  sg13g2_a22oi_1 _14807_ (
    .A1(_03260_),
    .A2(_04764_),
    .B1(_04766_),
    .B2(_04767_),
    .Y(_04768_)
  );
  sg13g2_o21ai_1 _14808_ (
    .A1(addr_i_5_),
    .A2(_00303_),
    .B1(addr_i_3_),
    .Y(_04769_)
  );
  sg13g2_o21ai_1 _14809_ (
    .A1(addr_i_3_),
    .A2(_02383_),
    .B1(_04769_),
    .Y(_04770_)
  );
  sg13g2_a221oi_1 _14810_ (
    .A1(addr_i_3_),
    .A2(_04139_),
    .B1(_04770_),
    .B2(_08011_),
    .C1(addr_i_7_),
    .Y(_04772_)
  );
  sg13g2_nor3_1 _14811_ (
    .A(_07293_),
    .B(_04768_),
    .C(_04772_),
    .Y(_04773_)
  );
  sg13g2_nor4_1 _14812_ (
    .A(_00243_),
    .B(_04758_),
    .C(_04763_),
    .D(_04773_),
    .Y(_04774_)
  );
  sg13g2_a22oi_1 _14813_ (
    .A1(_04736_),
    .A2(_04753_),
    .B1(_04774_),
    .B2(addr_i_10_),
    .Y(_04775_)
  );
  sg13g2_a21oi_1 _14814_ (
    .A1(_00476_),
    .A2(_01004_),
    .B1(_01520_),
    .Y(_04776_)
  );
  sg13g2_o21ai_1 _14815_ (
    .A1(_02419_),
    .A2(_04776_),
    .B1(_00061_),
    .Y(_04777_)
  );
  sg13g2_nor2_1 _14816_ (
    .A(_00016_),
    .B(_05678_),
    .Y(_04778_)
  );
  sg13g2_a21oi_1 _14817_ (
    .A1(_06873_),
    .A2(_01132_),
    .B1(_03260_),
    .Y(_04779_)
  );
  sg13g2_nor2_1 _14818_ (
    .A(_04778_),
    .B(_04779_),
    .Y(_04780_)
  );
  sg13g2_a21o_1 _14819_ (
    .A1(_04777_),
    .A2(_04780_),
    .B1(addr_i_6_),
    .X(_04781_)
  );
  sg13g2_or2_1 _14820_ (
    .A(_03186_),
    .B(_04130_),
    .X(_04783_)
  );
  sg13g2_a21oi_1 _14821_ (
    .A1(_00747_),
    .A2(_01144_),
    .B1(_03420_),
    .Y(_04784_)
  );
  sg13g2_a22oi_1 _14822_ (
    .A1(_09487_),
    .A2(_04783_),
    .B1(_04784_),
    .B2(addr_i_8_),
    .Y(_04785_)
  );
  sg13g2_nand2_1 _14823_ (
    .A(_00151_),
    .B(_00531_),
    .Y(_04786_)
  );
  sg13g2_a21o_1 _14824_ (
    .A1(addr_i_7_),
    .A2(_04786_),
    .B1(_02632_),
    .X(_04787_)
  );
  sg13g2_a21oi_1 _14825_ (
    .A1(_00403_),
    .A2(_07625_),
    .B1(_00961_),
    .Y(_04788_)
  );
  sg13g2_a21oi_1 _14826_ (
    .A1(_02369_),
    .A2(_01400_),
    .B1(_04788_),
    .Y(_04789_)
  );
  sg13g2_nor2_1 _14827_ (
    .A(addr_i_2_),
    .B(_04789_),
    .Y(_04790_)
  );
  sg13g2_o21ai_1 _14828_ (
    .A1(_00051_),
    .A2(_03229_),
    .B1(addr_i_8_),
    .Y(_04791_)
  );
  sg13g2_a22oi_1 _14829_ (
    .A1(_00827_),
    .A2(_04787_),
    .B1(_04790_),
    .B2(_04791_),
    .Y(_04792_)
  );
  sg13g2_a22oi_1 _14830_ (
    .A1(_04781_),
    .A2(_04785_),
    .B1(_04792_),
    .B2(_01211_),
    .Y(_04794_)
  );
  sg13g2_nor4_1 _14831_ (
    .A(addr_i_11_),
    .B(_04730_),
    .C(_04775_),
    .D(_04794_),
    .Y(_04795_)
  );
  sg13g2_nor2_1 _14832_ (
    .A(addr_i_7_),
    .B(_02033_),
    .Y(_04796_)
  );
  sg13g2_a21oi_1 _14833_ (
    .A1(_05645_),
    .A2(_01309_),
    .B1(_04796_),
    .Y(_04797_)
  );
  sg13g2_o21ai_1 _14834_ (
    .A1(_02040_),
    .A2(_04797_),
    .B1(addr_i_11_),
    .Y(_04798_)
  );
  sg13g2_nor2_1 _14835_ (
    .A(_09497_),
    .B(_00205_),
    .Y(_04799_)
  );
  sg13g2_o21ai_1 _14836_ (
    .A1(addr_i_3_),
    .A2(_04799_),
    .B1(_00567_),
    .Y(_04800_)
  );
  sg13g2_a21oi_1 _14837_ (
    .A1(_00704_),
    .A2(_02695_),
    .B1(_03260_),
    .Y(_04801_)
  );
  sg13g2_a22oi_1 _14838_ (
    .A1(_00123_),
    .A2(_04800_),
    .B1(_04801_),
    .B2(_01957_),
    .Y(_04802_)
  );
  sg13g2_nand2b_1 _14839_ (
    .A_N(_04802_),
    .B(_01119_),
    .Y(_04803_)
  );
  sg13g2_nand2_1 _14840_ (
    .A(_08388_),
    .B(_03458_),
    .Y(_04805_)
  );
  sg13g2_a21oi_1 _14841_ (
    .A1(_02187_),
    .A2(_04805_),
    .B1(addr_i_3_),
    .Y(_04806_)
  );
  sg13g2_a21o_1 _14842_ (
    .A1(_00607_),
    .A2(_01998_),
    .B1(_04806_),
    .X(_04807_)
  );
  sg13g2_o21ai_1 _14843_ (
    .A1(_03137_),
    .A2(_03565_),
    .B1(addr_i_3_),
    .Y(_04808_)
  );
  sg13g2_nand4_1 _14844_ (
    .A(_00223_),
    .B(_07625_),
    .C(_02513_),
    .D(_03226_),
    .Y(_04809_)
  );
  sg13g2_a21oi_1 _14845_ (
    .A1(_04808_),
    .A2(_04809_),
    .B1(_01034_),
    .Y(_04810_)
  );
  sg13g2_a22oi_1 _14846_ (
    .A1(_00277_),
    .A2(_04807_),
    .B1(_04810_),
    .B2(_01657_),
    .Y(_04811_)
  );
  sg13g2_xnor2_1 _14847_ (
    .A(_08774_),
    .B(_03466_),
    .Y(_04812_)
  );
  sg13g2_a221oi_1 _14848_ (
    .A1(_04803_),
    .A2(_04811_),
    .B1(_04812_),
    .B2(addr_i_9_),
    .C1(addr_i_10_),
    .Y(_04813_)
  );
  sg13g2_o21ai_1 _14849_ (
    .A1(_04798_),
    .A2(_04813_),
    .B1(addr_i_12_),
    .Y(_04814_)
  );
  sg13g2_a21oi_1 _14850_ (
    .A1(addr_i_3_),
    .A2(_02472_),
    .B1(_01881_),
    .Y(_04816_)
  );
  sg13g2_o21ai_1 _14851_ (
    .A1(_06717_),
    .A2(_04816_),
    .B1(_00430_),
    .Y(_04817_)
  );
  sg13g2_a21oi_1 _14852_ (
    .A1(addr_i_5_),
    .A2(_04817_),
    .B1(_04449_),
    .Y(_04818_)
  );
  sg13g2_nand2_1 _14853_ (
    .A(_01257_),
    .B(_00409_),
    .Y(_04819_)
  );
  sg13g2_a22oi_1 _14854_ (
    .A1(_02742_),
    .A2(_04819_),
    .B1(_02698_),
    .B2(addr_i_7_),
    .Y(_04820_)
  );
  sg13g2_nor2_1 _14855_ (
    .A(_04818_),
    .B(_04820_),
    .Y(_04821_)
  );
  sg13g2_o21ai_1 _14856_ (
    .A1(addr_i_3_),
    .A2(_03167_),
    .B1(_08520_),
    .Y(_04822_)
  );
  sg13g2_a21oi_1 _14857_ (
    .A1(addr_i_5_),
    .A2(_04822_),
    .B1(_03970_),
    .Y(_04823_)
  );
  sg13g2_o21ai_1 _14858_ (
    .A1(_08807_),
    .A2(_03153_),
    .B1(addr_i_4_),
    .Y(_04824_)
  );
  sg13g2_o21ai_1 _14859_ (
    .A1(addr_i_7_),
    .A2(_04823_),
    .B1(_04824_),
    .Y(_04825_)
  );
  sg13g2_nor2_1 _14860_ (
    .A(_09499_),
    .B(_00632_),
    .Y(_04827_)
  );
  sg13g2_a22oi_1 _14861_ (
    .A1(addr_i_7_),
    .A2(_03262_),
    .B1(_01231_),
    .B2(_03652_),
    .Y(_04828_)
  );
  sg13g2_a22oi_1 _14862_ (
    .A1(_01520_),
    .A2(_04827_),
    .B1(_04828_),
    .B2(_03260_),
    .Y(_04829_)
  );
  sg13g2_a21o_1 _14863_ (
    .A1(_02994_),
    .A2(_03882_),
    .B1(_00145_),
    .X(_04830_)
  );
  sg13g2_nor2_1 _14864_ (
    .A(addr_i_3_),
    .B(_04830_),
    .Y(_04831_)
  );
  sg13g2_a22oi_1 _14865_ (
    .A1(_00068_),
    .A2(_04825_),
    .B1(_04829_),
    .B2(_04831_),
    .Y(_04832_)
  );
  sg13g2_nor2_1 _14866_ (
    .A(_06706_),
    .B(_04832_),
    .Y(_04833_)
  );
  sg13g2_a22oi_1 _14867_ (
    .A1(_00114_),
    .A2(_04821_),
    .B1(_04833_),
    .B2(addr_i_9_),
    .Y(_04834_)
  );
  sg13g2_a21oi_1 _14868_ (
    .A1(addr_i_2_),
    .A2(_04572_),
    .B1(_09507_),
    .Y(_04835_)
  );
  sg13g2_a21oi_1 _14869_ (
    .A1(_01445_),
    .A2(_01231_),
    .B1(_00799_),
    .Y(_04836_)
  );
  sg13g2_o21ai_1 _14870_ (
    .A1(addr_i_4_),
    .A2(_04835_),
    .B1(_04836_),
    .Y(_04839_)
  );
  sg13g2_a221oi_1 _14871_ (
    .A1(_01159_),
    .A2(_00244_),
    .B1(_01215_),
    .B2(_00010_),
    .C1(addr_i_3_),
    .Y(_04840_)
  );
  sg13g2_inv_1 _14872_ (
    .A(_04840_),
    .Y(_04841_)
  );
  sg13g2_o21ai_1 _14873_ (
    .A1(_05292_),
    .A2(_02935_),
    .B1(_01131_),
    .Y(_04842_)
  );
  sg13g2_a21oi_1 _14874_ (
    .A1(_00651_),
    .A2(_04842_),
    .B1(_00324_),
    .Y(_04843_)
  );
  sg13g2_nor3_1 _14875_ (
    .A(addr_i_4_),
    .B(_00861_),
    .C(_01504_),
    .Y(_04844_)
  );
  sg13g2_nand2b_1 _14876_ (
    .A_N(_04844_),
    .B(addr_i_8_),
    .Y(_04845_)
  );
  sg13g2_a22oi_1 _14877_ (
    .A1(_04839_),
    .A2(_04841_),
    .B1(_04843_),
    .B2(_04845_),
    .Y(_04846_)
  );
  sg13g2_nor3_1 _14878_ (
    .A(_04108_),
    .B(addr_i_2_),
    .C(_03110_),
    .Y(_04847_)
  );
  sg13g2_a21oi_1 _14879_ (
    .A1(addr_i_2_),
    .A2(_00412_),
    .B1(_04847_),
    .Y(_04848_)
  );
  sg13g2_o21ai_1 _14880_ (
    .A1(_06795_),
    .A2(_09459_),
    .B1(_03690_),
    .Y(_04850_)
  );
  sg13g2_o21ai_1 _14881_ (
    .A1(_01615_),
    .A2(_04848_),
    .B1(_04850_),
    .Y(_04851_)
  );
  sg13g2_a21oi_1 _14882_ (
    .A1(_09510_),
    .A2(_06784_),
    .B1(addr_i_2_),
    .Y(_04852_)
  );
  sg13g2_nor2_1 _14883_ (
    .A(_00946_),
    .B(_04852_),
    .Y(_04853_)
  );
  sg13g2_nand2_1 _14884_ (
    .A(_02089_),
    .B(_01004_),
    .Y(_04854_)
  );
  sg13g2_nor2_1 _14885_ (
    .A(addr_i_4_),
    .B(_04854_),
    .Y(_04855_)
  );
  sg13g2_a22oi_1 _14886_ (
    .A1(addr_i_4_),
    .A2(_04853_),
    .B1(_04855_),
    .B2(addr_i_3_),
    .Y(_04856_)
  );
  sg13g2_nand2_1 _14887_ (
    .A(_00113_),
    .B(_02149_),
    .Y(_04857_)
  );
  sg13g2_a22oi_1 _14888_ (
    .A1(addr_i_3_),
    .A2(_04851_),
    .B1(_04856_),
    .B2(_04857_),
    .Y(_04858_)
  );
  sg13g2_o21ai_1 _14889_ (
    .A1(_04846_),
    .A2(_04858_),
    .B1(addr_i_9_),
    .Y(_04859_)
  );
  sg13g2_nand2_1 _14890_ (
    .A(_00511_),
    .B(_04859_),
    .Y(_04861_)
  );
  sg13g2_nor2_1 _14891_ (
    .A(_04108_),
    .B(_07061_),
    .Y(_04862_)
  );
  sg13g2_o21ai_1 _14892_ (
    .A1(_03914_),
    .A2(_04862_),
    .B1(_06154_),
    .Y(_04863_)
  );
  sg13g2_nor3_1 _14893_ (
    .A(_00115_),
    .B(_05568_),
    .C(_00632_),
    .Y(_04864_)
  );
  sg13g2_a22oi_1 _14894_ (
    .A1(_00701_),
    .A2(_04863_),
    .B1(_04864_),
    .B2(addr_i_6_),
    .Y(_04865_)
  );
  sg13g2_nand2_1 _14895_ (
    .A(_03665_),
    .B(_01570_),
    .Y(_04866_)
  );
  sg13g2_a21o_1 _14896_ (
    .A1(_00566_),
    .A2(_04866_),
    .B1(addr_i_2_),
    .X(_04867_)
  );
  sg13g2_a21oi_1 _14897_ (
    .A1(_01708_),
    .A2(_04867_),
    .B1(addr_i_7_),
    .Y(_04868_)
  );
  sg13g2_a22oi_1 _14898_ (
    .A1(_00169_),
    .A2(_00177_),
    .B1(_04865_),
    .B2(_04868_),
    .Y(_04869_)
  );
  sg13g2_a22oi_1 _14899_ (
    .A1(_01881_),
    .A2(_07038_),
    .B1(_02639_),
    .B2(addr_i_5_),
    .Y(_04870_)
  );
  sg13g2_a221oi_1 _14900_ (
    .A1(_09492_),
    .A2(_00616_),
    .B1(_04720_),
    .B2(addr_i_3_),
    .C1(_02063_),
    .Y(_04872_)
  );
  sg13g2_o21ai_1 _14901_ (
    .A1(_04870_),
    .A2(_04872_),
    .B1(addr_i_2_),
    .Y(_04873_)
  );
  sg13g2_and2_1 _14902_ (
    .A(_01008_),
    .B(_01734_),
    .X(_04874_)
  );
  sg13g2_a22oi_1 _14903_ (
    .A1(_00428_),
    .A2(_03348_),
    .B1(_03880_),
    .B2(addr_i_2_),
    .Y(_04875_)
  );
  sg13g2_o21ai_1 _14904_ (
    .A1(addr_i_3_),
    .A2(_04874_),
    .B1(_04875_),
    .Y(_04876_)
  );
  sg13g2_a21oi_1 _14905_ (
    .A1(_04873_),
    .A2(_04876_),
    .B1(_07293_),
    .Y(_04877_)
  );
  sg13g2_a21oi_1 _14906_ (
    .A1(_06706_),
    .A2(_04869_),
    .B1(_04877_),
    .Y(_04878_)
  );
  sg13g2_o21ai_1 _14907_ (
    .A1(addr_i_4_),
    .A2(_01789_),
    .B1(_00651_),
    .Y(_04879_)
  );
  sg13g2_a22oi_1 _14908_ (
    .A1(_05877_),
    .A2(_04879_),
    .B1(_00518_),
    .B2(_00290_),
    .Y(_04880_)
  );
  sg13g2_nand2_1 _14909_ (
    .A(_04528_),
    .B(_05225_),
    .Y(_04881_)
  );
  sg13g2_nand3_1 _14910_ (
    .A(_00150_),
    .B(_01301_),
    .C(_00386_),
    .Y(_04883_)
  );
  sg13g2_nand2_1 _14911_ (
    .A(_04881_),
    .B(_04883_),
    .Y(_04884_)
  );
  sg13g2_a21oi_1 _14912_ (
    .A1(_01203_),
    .A2(_02738_),
    .B1(addr_i_3_),
    .Y(_04885_)
  );
  sg13g2_o21ai_1 _14913_ (
    .A1(_02238_),
    .A2(_00977_),
    .B1(_00305_),
    .Y(_04886_)
  );
  sg13g2_nand3_1 _14914_ (
    .A(_06695_),
    .B(_00980_),
    .C(_04886_),
    .Y(_04887_)
  );
  sg13g2_a22oi_1 _14915_ (
    .A1(addr_i_3_),
    .A2(_04884_),
    .B1(_04885_),
    .B2(_04887_),
    .Y(_04888_)
  );
  sg13g2_nand3b_1 _14916_ (
    .A_N(_04757_),
    .B(addr_i_4_),
    .C(_00211_),
    .Y(_04889_)
  );
  sg13g2_nand3_1 _14917_ (
    .A(_01095_),
    .B(_03575_),
    .C(_02077_),
    .Y(_04890_)
  );
  sg13g2_a21oi_1 _14918_ (
    .A1(_04889_),
    .A2(_04890_),
    .B1(_08487_),
    .Y(_04891_)
  );
  sg13g2_nor4_1 _14919_ (
    .A(_00925_),
    .B(_04880_),
    .C(_04888_),
    .D(_04891_),
    .Y(_04892_)
  );
  sg13g2_a22oi_1 _14920_ (
    .A1(_01176_),
    .A2(_04878_),
    .B1(_04892_),
    .B2(addr_i_11_),
    .Y(_04894_)
  );
  sg13g2_o21ai_1 _14921_ (
    .A1(_04834_),
    .A2(_04861_),
    .B1(_04894_),
    .Y(_04895_)
  );
  sg13g2_o21ai_1 _14922_ (
    .A1(_06419_),
    .A2(_00010_),
    .B1(_00951_),
    .Y(_04896_)
  );
  sg13g2_a21oi_1 _14923_ (
    .A1(_09513_),
    .A2(_02319_),
    .B1(addr_i_5_),
    .Y(_04897_)
  );
  sg13g2_a21oi_1 _14924_ (
    .A1(_00401_),
    .A2(_04896_),
    .B1(_04897_),
    .Y(_04898_)
  );
  sg13g2_o21ai_1 _14925_ (
    .A1(_00467_),
    .A2(_02437_),
    .B1(_04898_),
    .Y(_04899_)
  );
  sg13g2_a21oi_1 _14926_ (
    .A1(_04162_),
    .A2(_08930_),
    .B1(_04461_),
    .Y(_04900_)
  );
  sg13g2_o21ai_1 _14927_ (
    .A1(_00474_),
    .A2(_04900_),
    .B1(addr_i_4_),
    .Y(_04901_)
  );
  sg13g2_a21oi_1 _14928_ (
    .A1(_00131_),
    .A2(_04901_),
    .B1(addr_i_7_),
    .Y(_04902_)
  );
  sg13g2_o21ai_1 _14929_ (
    .A1(_08553_),
    .A2(_00973_),
    .B1(addr_i_8_),
    .Y(_04903_)
  );
  sg13g2_a22oi_1 _14930_ (
    .A1(addr_i_2_),
    .A2(_04899_),
    .B1(_04902_),
    .B2(_04903_),
    .Y(_04905_)
  );
  sg13g2_nor3_1 _14931_ (
    .A(addr_i_4_),
    .B(addr_i_2_),
    .C(_00011_),
    .Y(_04906_)
  );
  sg13g2_nor2_1 _14932_ (
    .A(_01277_),
    .B(_04906_),
    .Y(_04907_)
  );
  sg13g2_nand2_1 _14933_ (
    .A(_04164_),
    .B(_04907_),
    .Y(_04908_)
  );
  sg13g2_nor2_1 _14934_ (
    .A(_01212_),
    .B(_03478_),
    .Y(_04909_)
  );
  sg13g2_a22oi_1 _14935_ (
    .A1(_01475_),
    .A2(_04908_),
    .B1(_04909_),
    .B2(_00191_),
    .Y(_04910_)
  );
  sg13g2_o21ai_1 _14936_ (
    .A1(_07337_),
    .A2(_05247_),
    .B1(_01729_),
    .Y(_04911_)
  );
  sg13g2_a221oi_1 _14937_ (
    .A1(_03690_),
    .A2(_00745_),
    .B1(_04911_),
    .B2(addr_i_4_),
    .C1(addr_i_3_),
    .Y(_04912_)
  );
  sg13g2_o21ai_1 _14938_ (
    .A1(_04910_),
    .A2(_04912_),
    .B1(_02576_),
    .Y(_04913_)
  );
  sg13g2_nand3b_1 _14939_ (
    .A_N(_04905_),
    .B(_05214_),
    .C(_04913_),
    .Y(_04914_)
  );
  sg13g2_nand2_1 _14940_ (
    .A(_06054_),
    .B(_06099_),
    .Y(_04916_)
  );
  sg13g2_o21ai_1 _14941_ (
    .A1(_04139_),
    .A2(_04906_),
    .B1(addr_i_3_),
    .Y(_04917_)
  );
  sg13g2_a21oi_1 _14942_ (
    .A1(_06862_),
    .A2(_02683_),
    .B1(addr_i_3_),
    .Y(_04918_)
  );
  sg13g2_o21ai_1 _14943_ (
    .A1(_03577_),
    .A2(_04918_),
    .B1(addr_i_5_),
    .Y(_04919_)
  );
  sg13g2_nand3_1 _14944_ (
    .A(_04916_),
    .B(_04917_),
    .C(_04919_),
    .Y(_04920_)
  );
  sg13g2_nand3_1 _14945_ (
    .A(_01878_),
    .B(_09479_),
    .C(_00832_),
    .Y(_04921_)
  );
  sg13g2_a21oi_1 _14946_ (
    .A1(_00650_),
    .A2(_09475_),
    .B1(addr_i_3_),
    .Y(_04922_)
  );
  sg13g2_o21ai_1 _14947_ (
    .A1(_02922_),
    .A2(_04922_),
    .B1(_05247_),
    .Y(_04923_)
  );
  sg13g2_nand3_1 _14948_ (
    .A(addr_i_8_),
    .B(_04921_),
    .C(_04923_),
    .Y(_04924_)
  );
  sg13g2_a21oi_1 _14949_ (
    .A1(addr_i_7_),
    .A2(_04920_),
    .B1(_04924_),
    .Y(_04925_)
  );
  sg13g2_a21oi_1 _14950_ (
    .A1(_00032_),
    .A2(_01704_),
    .B1(addr_i_5_),
    .Y(_04927_)
  );
  sg13g2_nor2_1 _14951_ (
    .A(_01686_),
    .B(_04927_),
    .Y(_04928_)
  );
  sg13g2_a21oi_1 _14952_ (
    .A1(_00047_),
    .A2(_04874_),
    .B1(_04928_),
    .Y(_04929_)
  );
  sg13g2_a21oi_1 _14953_ (
    .A1(_03993_),
    .A2(_00301_),
    .B1(_00029_),
    .Y(_04930_)
  );
  sg13g2_a21oi_1 _14954_ (
    .A1(_03993_),
    .A2(_00029_),
    .B1(addr_i_8_),
    .Y(_04931_)
  );
  sg13g2_o21ai_1 _14955_ (
    .A1(addr_i_4_),
    .A2(_04930_),
    .B1(_04931_),
    .Y(_04932_)
  );
  sg13g2_nand2_1 _14956_ (
    .A(addr_i_3_),
    .B(_01539_),
    .Y(_04933_)
  );
  sg13g2_o21ai_1 _14957_ (
    .A1(_08056_),
    .A2(_03033_),
    .B1(addr_i_2_),
    .Y(_04934_)
  );
  sg13g2_a21oi_1 _14958_ (
    .A1(_04933_),
    .A2(_04934_),
    .B1(_00053_),
    .Y(_04935_)
  );
  sg13g2_a22oi_1 _14959_ (
    .A1(addr_i_2_),
    .A2(_04929_),
    .B1(_04932_),
    .B2(_04935_),
    .Y(_04936_)
  );
  sg13g2_or3_1 _14960_ (
    .A(_06652_),
    .B(_04925_),
    .C(_04936_),
    .X(_04938_)
  );
  sg13g2_a21oi_1 _14961_ (
    .A1(_02250_),
    .A2(_01084_),
    .B1(addr_i_3_),
    .Y(_04939_)
  );
  sg13g2_o21ai_1 _14962_ (
    .A1(_01202_),
    .A2(_04939_),
    .B1(_02501_),
    .Y(_04940_)
  );
  sg13g2_nor2_1 _14963_ (
    .A(_01292_),
    .B(_07193_),
    .Y(_04941_)
  );
  sg13g2_o21ai_1 _14964_ (
    .A1(addr_i_3_),
    .A2(_04941_),
    .B1(addr_i_8_),
    .Y(_04942_)
  );
  sg13g2_nand2_1 _14965_ (
    .A(_00242_),
    .B(_00210_),
    .Y(_04943_)
  );
  sg13g2_a21oi_1 _14966_ (
    .A1(_00846_),
    .A2(_04943_),
    .B1(_02277_),
    .Y(_04944_)
  );
  sg13g2_o21ai_1 _14967_ (
    .A1(_01202_),
    .A2(_00649_),
    .B1(addr_i_6_),
    .Y(_04945_)
  );
  sg13g2_a22oi_1 _14968_ (
    .A1(addr_i_3_),
    .A2(_00338_),
    .B1(_02055_),
    .B2(addr_i_8_),
    .Y(_04946_)
  );
  sg13g2_a21oi_1 _14969_ (
    .A1(_04945_),
    .A2(_04946_),
    .B1(addr_i_7_),
    .Y(_04947_)
  );
  sg13g2_o21ai_1 _14970_ (
    .A1(_04942_),
    .A2(_04944_),
    .B1(_04947_),
    .Y(_04950_)
  );
  sg13g2_o21ai_1 _14971_ (
    .A1(_02479_),
    .A2(_02498_),
    .B1(_01160_),
    .Y(_04951_)
  );
  sg13g2_nor2_1 _14972_ (
    .A(addr_i_5_),
    .B(_01914_),
    .Y(_04952_)
  );
  sg13g2_a22oi_1 _14973_ (
    .A1(addr_i_3_),
    .A2(_04951_),
    .B1(_04952_),
    .B2(_00825_),
    .Y(_04953_)
  );
  sg13g2_a21oi_1 _14974_ (
    .A1(addr_i_5_),
    .A2(_02498_),
    .B1(_00692_),
    .Y(_04954_)
  );
  sg13g2_o21ai_1 _14975_ (
    .A1(_00491_),
    .A2(_04954_),
    .B1(addr_i_4_),
    .Y(_04955_)
  );
  sg13g2_nand2_1 _14976_ (
    .A(_04953_),
    .B(_04955_),
    .Y(_04956_)
  );
  sg13g2_a21oi_1 _14977_ (
    .A1(addr_i_2_),
    .A2(_02722_),
    .B1(addr_i_5_),
    .Y(_04957_)
  );
  sg13g2_o21ai_1 _14978_ (
    .A1(_02923_),
    .A2(_04957_),
    .B1(_01047_),
    .Y(_04958_)
  );
  sg13g2_nand4_1 _14979_ (
    .A(_04940_),
    .B(_04950_),
    .C(_04956_),
    .D(_04958_),
    .Y(_04959_)
  );
  sg13g2_nor2_1 _14980_ (
    .A(_01656_),
    .B(_00951_),
    .Y(_04961_)
  );
  sg13g2_nand3_1 _14981_ (
    .A(addr_i_3_),
    .B(_01672_),
    .C(_00284_),
    .Y(_04962_)
  );
  sg13g2_a21oi_1 _14982_ (
    .A1(_01945_),
    .A2(_04962_),
    .B1(_09271_),
    .Y(_04963_)
  );
  sg13g2_o21ai_1 _14983_ (
    .A1(_04961_),
    .A2(_04963_),
    .B1(addr_i_5_),
    .Y(_04964_)
  );
  sg13g2_o21ai_1 _14984_ (
    .A1(_00959_),
    .A2(_00110_),
    .B1(addr_i_6_),
    .Y(_04965_)
  );
  sg13g2_nor3_1 _14985_ (
    .A(_04981_),
    .B(_03577_),
    .C(_00247_),
    .Y(_04966_)
  );
  sg13g2_a22oi_1 _14986_ (
    .A1(_00910_),
    .A2(_04965_),
    .B1(_04966_),
    .B2(addr_i_5_),
    .Y(_04967_)
  );
  sg13g2_a22oi_1 _14987_ (
    .A1(_00073_),
    .A2(_00100_),
    .B1(_01611_),
    .B2(_04967_),
    .Y(_04968_)
  );
  sg13g2_nand2_1 _14988_ (
    .A(_00347_),
    .B(_01097_),
    .Y(_04969_)
  );
  sg13g2_o21ai_1 _14989_ (
    .A1(addr_i_2_),
    .A2(_01304_),
    .B1(_04969_),
    .Y(_04970_)
  );
  sg13g2_o21ai_1 _14990_ (
    .A1(_00007_),
    .A2(_00105_),
    .B1(_00422_),
    .Y(_04972_)
  );
  sg13g2_nor4_1 _14991_ (
    .A(_01155_),
    .B(_00503_),
    .C(_00569_),
    .D(_02850_),
    .Y(_04973_)
  );
  sg13g2_a22oi_1 _14992_ (
    .A1(_01320_),
    .A2(_04970_),
    .B1(_04972_),
    .B2(_04973_),
    .Y(_04974_)
  );
  sg13g2_nor2_1 _14993_ (
    .A(_00060_),
    .B(_02241_),
    .Y(_04975_)
  );
  sg13g2_o21ai_1 _14994_ (
    .A1(_01846_),
    .A2(_04975_),
    .B1(_00402_),
    .Y(_04976_)
  );
  sg13g2_a221oi_1 _14995_ (
    .A1(_04964_),
    .A2(_04968_),
    .B1(_04974_),
    .B2(_04976_),
    .C1(addr_i_10_),
    .Y(_04977_)
  );
  sg13g2_o21ai_1 _14996_ (
    .A1(_00397_),
    .A2(_04959_),
    .B1(_04977_),
    .Y(_04978_)
  );
  sg13g2_nand4_1 _14997_ (
    .A(addr_i_11_),
    .B(_04914_),
    .C(_04938_),
    .D(_04978_),
    .Y(_04979_)
  );
  sg13g2_nand3_1 _14998_ (
    .A(_02251_),
    .B(_04895_),
    .C(_04979_),
    .Y(_04980_)
  );
  sg13g2_o21ai_1 _14999_ (
    .A1(_04795_),
    .A2(_04814_),
    .B1(_04980_),
    .Y(data_o_22_)
  );
  sg13g2_a21oi_1 _15000_ (
    .A1(_02213_),
    .A2(_01791_),
    .B1(_00145_),
    .Y(_04982_)
  );
  sg13g2_nor2_1 _15001_ (
    .A(_03152_),
    .B(_04982_),
    .Y(_04983_)
  );
  sg13g2_a22oi_1 _15002_ (
    .A1(addr_i_2_),
    .A2(_01154_),
    .B1(_02198_),
    .B2(addr_i_4_),
    .Y(_04984_)
  );
  sg13g2_a22oi_1 _15003_ (
    .A1(addr_i_4_),
    .A2(_04983_),
    .B1(_04984_),
    .B2(_05877_),
    .Y(_04985_)
  );
  sg13g2_nand2_1 _15004_ (
    .A(_00351_),
    .B(_05081_),
    .Y(_04986_)
  );
  sg13g2_o21ai_1 _15005_ (
    .A1(_01567_),
    .A2(_03382_),
    .B1(_04191_),
    .Y(_04987_)
  );
  sg13g2_a21oi_1 _15006_ (
    .A1(_04986_),
    .A2(_04987_),
    .B1(addr_i_3_),
    .Y(_04988_)
  );
  sg13g2_a22oi_1 _15007_ (
    .A1(_00500_),
    .A2(_00029_),
    .B1(_04985_),
    .B2(_04988_),
    .Y(_04989_)
  );
  sg13g2_nand2b_1 _15008_ (
    .A_N(_04989_),
    .B(addr_i_8_),
    .Y(_04990_)
  );
  sg13g2_nand3_1 _15009_ (
    .A(_00360_),
    .B(_07337_),
    .C(_01367_),
    .Y(_04991_)
  );
  sg13g2_nand2_1 _15010_ (
    .A(_02472_),
    .B(_02732_),
    .Y(_04993_)
  );
  sg13g2_nor2_1 _15011_ (
    .A(_01615_),
    .B(_04993_),
    .Y(_04994_)
  );
  sg13g2_a22oi_1 _15012_ (
    .A1(_01413_),
    .A2(_04991_),
    .B1(_04994_),
    .B2(_05877_),
    .Y(_04995_)
  );
  sg13g2_a21o_1 _15013_ (
    .A1(addr_i_5_),
    .A2(_01264_),
    .B1(_00818_),
    .X(_04996_)
  );
  sg13g2_nor2_1 _15014_ (
    .A(_01815_),
    .B(_01486_),
    .Y(_04997_)
  );
  sg13g2_a22oi_1 _15015_ (
    .A1(addr_i_7_),
    .A2(_04996_),
    .B1(_04997_),
    .B2(addr_i_3_),
    .Y(_04998_)
  );
  sg13g2_or4_1 _15016_ (
    .A(addr_i_8_),
    .B(_04499_),
    .C(_04995_),
    .D(_04998_),
    .X(_04999_)
  );
  sg13g2_a21oi_1 _15017_ (
    .A1(_04990_),
    .A2(_04999_),
    .B1(_00109_),
    .Y(_05000_)
  );
  sg13g2_a21oi_1 _15018_ (
    .A1(addr_i_4_),
    .A2(_07326_),
    .B1(addr_i_6_),
    .Y(_05001_)
  );
  sg13g2_a21oi_1 _15019_ (
    .A1(_00731_),
    .A2(_00571_),
    .B1(addr_i_5_),
    .Y(_05002_)
  );
  sg13g2_a22oi_1 _15020_ (
    .A1(addr_i_3_),
    .A2(_01815_),
    .B1(_05001_),
    .B2(_05002_),
    .Y(_05004_)
  );
  sg13g2_and2_1 _15021_ (
    .A(_04119_),
    .B(_06983_),
    .X(_05005_)
  );
  sg13g2_o21ai_1 _15022_ (
    .A1(_03587_),
    .A2(_05005_),
    .B1(_06375_),
    .Y(_05006_)
  );
  sg13g2_o21ai_1 _15023_ (
    .A1(_01615_),
    .A2(_05004_),
    .B1(_05006_),
    .Y(_05007_)
  );
  sg13g2_a21oi_1 _15024_ (
    .A1(_01527_),
    .A2(_08022_),
    .B1(addr_i_6_),
    .Y(_05008_)
  );
  sg13g2_a21oi_1 _15025_ (
    .A1(_00156_),
    .A2(_00917_),
    .B1(_05008_),
    .Y(_05009_)
  );
  sg13g2_nor3_1 _15026_ (
    .A(addr_i_4_),
    .B(_07812_),
    .C(_07636_),
    .Y(_05010_)
  );
  sg13g2_a22oi_1 _15027_ (
    .A1(addr_i_3_),
    .A2(_02057_),
    .B1(_05010_),
    .B2(_00791_),
    .Y(_05011_)
  );
  sg13g2_o21ai_1 _15028_ (
    .A1(addr_i_6_),
    .A2(_05335_),
    .B1(addr_i_4_),
    .Y(_05012_)
  );
  sg13g2_nor2_1 _15029_ (
    .A(_01276_),
    .B(_02423_),
    .Y(_05013_)
  );
  sg13g2_a21o_1 _15030_ (
    .A1(_05012_),
    .A2(_05013_),
    .B1(addr_i_3_),
    .X(_05015_)
  );
  sg13g2_nor2_1 _15031_ (
    .A(_02424_),
    .B(_01244_),
    .Y(_05016_)
  );
  sg13g2_a21oi_1 _15032_ (
    .A1(_00039_),
    .A2(_05016_),
    .B1(_08045_),
    .Y(_05017_)
  );
  sg13g2_a21oi_1 _15033_ (
    .A1(_05011_),
    .A2(_05015_),
    .B1(_05017_),
    .Y(_05018_)
  );
  sg13g2_o21ai_1 _15034_ (
    .A1(_00860_),
    .A2(_05009_),
    .B1(_05018_),
    .Y(_05019_)
  );
  sg13g2_a21o_1 _15035_ (
    .A1(addr_i_8_),
    .A2(_05007_),
    .B1(_05019_),
    .X(_05020_)
  );
  sg13g2_nor2_1 _15036_ (
    .A(_00342_),
    .B(_00676_),
    .Y(_05021_)
  );
  sg13g2_o21ai_1 _15037_ (
    .A1(addr_i_2_),
    .A2(_05021_),
    .B1(_02528_),
    .Y(_05022_)
  );
  sg13g2_nand3_1 _15038_ (
    .A(addr_i_3_),
    .B(_02694_),
    .C(_02467_),
    .Y(_05023_)
  );
  sg13g2_o21ai_1 _15039_ (
    .A1(addr_i_3_),
    .A2(_05022_),
    .B1(_05023_),
    .Y(_05024_)
  );
  sg13g2_nand3_1 _15040_ (
    .A(addr_i_4_),
    .B(_00703_),
    .C(_00747_),
    .Y(_05026_)
  );
  sg13g2_a21oi_1 _15041_ (
    .A1(_05024_),
    .A2(_05026_),
    .B1(_02535_),
    .Y(_05027_)
  );
  sg13g2_nor3_1 _15042_ (
    .A(_00128_),
    .B(_04062_),
    .C(_04906_),
    .Y(_05028_)
  );
  sg13g2_a21oi_1 _15043_ (
    .A1(_01125_),
    .A2(_03457_),
    .B1(_00967_),
    .Y(_05029_)
  );
  sg13g2_a22oi_1 _15044_ (
    .A1(_04442_),
    .A2(_01179_),
    .B1(_03494_),
    .B2(_05029_),
    .Y(_05030_)
  );
  sg13g2_o21ai_1 _15045_ (
    .A1(addr_i_3_),
    .A2(_05028_),
    .B1(_05030_),
    .Y(_05031_)
  );
  sg13g2_o21ai_1 _15046_ (
    .A1(_00159_),
    .A2(_02374_),
    .B1(_02530_),
    .Y(_05032_)
  );
  sg13g2_o21ai_1 _15047_ (
    .A1(_01282_),
    .A2(_00569_),
    .B1(addr_i_6_),
    .Y(_05033_)
  );
  sg13g2_a22oi_1 _15048_ (
    .A1(_01519_),
    .A2(_01830_),
    .B1(_02963_),
    .B2(_00227_),
    .Y(_05034_)
  );
  sg13g2_nand3_1 _15049_ (
    .A(_05032_),
    .B(_05033_),
    .C(_05034_),
    .Y(_05035_)
  );
  sg13g2_nor2_1 _15050_ (
    .A(addr_i_5_),
    .B(_05524_),
    .Y(_05037_)
  );
  sg13g2_nor2_1 _15051_ (
    .A(_02990_),
    .B(_05037_),
    .Y(_05038_)
  );
  sg13g2_o21ai_1 _15052_ (
    .A1(_00015_),
    .A2(_05038_),
    .B1(addr_i_6_),
    .Y(_05039_)
  );
  sg13g2_o21ai_1 _15053_ (
    .A1(_00626_),
    .A2(_00947_),
    .B1(addr_i_4_),
    .Y(_05040_)
  );
  sg13g2_nand4_1 _15054_ (
    .A(_00148_),
    .B(_03890_),
    .C(_05039_),
    .D(_05040_),
    .Y(_05041_)
  );
  sg13g2_nand3_1 _15055_ (
    .A(_05031_),
    .B(_05035_),
    .C(_05041_),
    .Y(_05042_)
  );
  sg13g2_a22oi_1 _15056_ (
    .A1(addr_i_9_),
    .A2(_05020_),
    .B1(_05027_),
    .B2(_05042_),
    .Y(_05043_)
  );
  sg13g2_a21oi_1 _15057_ (
    .A1(addr_i_7_),
    .A2(_00749_),
    .B1(addr_i_5_),
    .Y(_05044_)
  );
  sg13g2_a22oi_1 _15058_ (
    .A1(addr_i_3_),
    .A2(_03723_),
    .B1(_05044_),
    .B2(_09507_),
    .Y(_05045_)
  );
  sg13g2_nand2_1 _15059_ (
    .A(_01738_),
    .B(_00620_),
    .Y(_05046_)
  );
  sg13g2_o21ai_1 _15060_ (
    .A1(addr_i_5_),
    .A2(_07105_),
    .B1(addr_i_2_),
    .Y(_05048_)
  );
  sg13g2_a21oi_1 _15061_ (
    .A1(_00520_),
    .A2(_05048_),
    .B1(addr_i_3_),
    .Y(_05049_)
  );
  sg13g2_o21ai_1 _15062_ (
    .A1(_02064_),
    .A2(_01628_),
    .B1(_09260_),
    .Y(_05050_)
  );
  sg13g2_a22oi_1 _15063_ (
    .A1(addr_i_3_),
    .A2(_05046_),
    .B1(_05049_),
    .B2(_05050_),
    .Y(_05051_)
  );
  sg13g2_mux2_1 _15064_ (
    .A0(_05045_),
    .A1(_05051_),
    .S(addr_i_4_),
    .X(_05052_)
  );
  sg13g2_a22oi_1 _15065_ (
    .A1(_01282_),
    .A2(_09487_),
    .B1(_00632_),
    .B2(addr_i_8_),
    .Y(_05053_)
  );
  sg13g2_o21ai_1 _15066_ (
    .A1(_02154_),
    .A2(_04276_),
    .B1(addr_i_3_),
    .Y(_05054_)
  );
  sg13g2_nand3_1 _15067_ (
    .A(_00146_),
    .B(_03391_),
    .C(_05054_),
    .Y(_05055_)
  );
  sg13g2_o21ai_1 _15068_ (
    .A1(addr_i_6_),
    .A2(_01587_),
    .B1(_00156_),
    .Y(_05056_)
  );
  sg13g2_o21ai_1 _15069_ (
    .A1(_00838_),
    .A2(_02514_),
    .B1(addr_i_7_),
    .Y(_05057_)
  );
  sg13g2_nand2_1 _15070_ (
    .A(_00799_),
    .B(_03152_),
    .Y(_05060_)
  );
  sg13g2_nand4_1 _15071_ (
    .A(addr_i_2_),
    .B(_05056_),
    .C(_05057_),
    .D(_05060_),
    .Y(_05061_)
  );
  sg13g2_nor2_1 _15072_ (
    .A(addr_i_3_),
    .B(_03112_),
    .Y(_05062_)
  );
  sg13g2_o21ai_1 _15073_ (
    .A1(_01543_),
    .A2(_00594_),
    .B1(_03652_),
    .Y(_05063_)
  );
  sg13g2_a21oi_1 _15074_ (
    .A1(_01948_),
    .A2(_00764_),
    .B1(_00565_),
    .Y(_05064_)
  );
  sg13g2_nor3_1 _15075_ (
    .A(_05062_),
    .B(_05063_),
    .C(_05064_),
    .Y(_05065_)
  );
  sg13g2_o21ai_1 _15076_ (
    .A1(_00185_),
    .A2(_03497_),
    .B1(addr_i_8_),
    .Y(_05066_)
  );
  sg13g2_a22oi_1 _15077_ (
    .A1(_05055_),
    .A2(_05061_),
    .B1(_05065_),
    .B2(_05066_),
    .Y(_05067_)
  );
  sg13g2_a22oi_1 _15078_ (
    .A1(_05052_),
    .A2(_05053_),
    .B1(_06652_),
    .B2(_05067_),
    .Y(_05068_)
  );
  sg13g2_nor2_1 _15079_ (
    .A(addr_i_11_),
    .B(_05068_),
    .Y(_05069_)
  );
  sg13g2_o21ai_1 _15080_ (
    .A1(addr_i_10_),
    .A2(_05043_),
    .B1(_05069_),
    .Y(_05071_)
  );
  sg13g2_nor2_1 _15081_ (
    .A(_06684_),
    .B(_01159_),
    .Y(_05072_)
  );
  sg13g2_xnor2_1 _15082_ (
    .A(_00701_),
    .B(_05072_),
    .Y(_05073_)
  );
  sg13g2_a21oi_1 _15083_ (
    .A1(addr_i_9_),
    .A2(_05073_),
    .B1(addr_i_10_),
    .Y(_05074_)
  );
  sg13g2_o21ai_1 _15084_ (
    .A1(_00156_),
    .A2(_00474_),
    .B1(addr_i_2_),
    .Y(_05075_)
  );
  sg13g2_nand2_1 _15085_ (
    .A(_00371_),
    .B(_02634_),
    .Y(_05076_)
  );
  sg13g2_a21oi_1 _15086_ (
    .A1(addr_i_3_),
    .A2(_05076_),
    .B1(_05932_),
    .Y(_05077_)
  );
  sg13g2_nand3_1 _15087_ (
    .A(_02434_),
    .B(_05075_),
    .C(_05077_),
    .Y(_05078_)
  );
  sg13g2_nand2_1 _15088_ (
    .A(_00688_),
    .B(_01398_),
    .Y(_05079_)
  );
  sg13g2_a22oi_1 _15089_ (
    .A1(addr_i_2_),
    .A2(_05079_),
    .B1(_00009_),
    .B2(_01481_),
    .Y(_05080_)
  );
  sg13g2_a22oi_1 _15090_ (
    .A1(addr_i_7_),
    .A2(_05078_),
    .B1(_05080_),
    .B2(addr_i_8_),
    .Y(_05082_)
  );
  sg13g2_nand2_1 _15091_ (
    .A(_04119_),
    .B(_09485_),
    .Y(_05083_)
  );
  sg13g2_nand2_1 _15092_ (
    .A(_01709_),
    .B(_05083_),
    .Y(_05084_)
  );
  sg13g2_nor3_1 _15093_ (
    .A(addr_i_6_),
    .B(_04539_),
    .C(_00951_),
    .Y(_05085_)
  );
  sg13g2_a21o_1 _15094_ (
    .A1(addr_i_4_),
    .A2(_05084_),
    .B1(_05085_),
    .X(_05086_)
  );
  sg13g2_nand3_1 _15095_ (
    .A(_02063_),
    .B(_02472_),
    .C(_00155_),
    .Y(_05087_)
  );
  sg13g2_nand3_1 _15096_ (
    .A(_05822_),
    .B(_02467_),
    .C(_05087_),
    .Y(_05088_)
  );
  sg13g2_o21ai_1 _15097_ (
    .A1(_08011_),
    .A2(_02987_),
    .B1(addr_i_8_),
    .Y(_05089_)
  );
  sg13g2_a221oi_1 _15098_ (
    .A1(addr_i_5_),
    .A2(_05086_),
    .B1(_05088_),
    .B2(addr_i_3_),
    .C1(_05089_),
    .Y(_05090_)
  );
  sg13g2_o21ai_1 _15099_ (
    .A1(_06795_),
    .A2(_00617_),
    .B1(addr_i_3_),
    .Y(_05091_)
  );
  sg13g2_nand3_1 _15100_ (
    .A(_00224_),
    .B(_01378_),
    .C(_05091_),
    .Y(_05093_)
  );
  sg13g2_and2_1 _15101_ (
    .A(_02700_),
    .B(_05093_),
    .X(_05094_)
  );
  sg13g2_o21ai_1 _15102_ (
    .A1(_05082_),
    .A2(_05090_),
    .B1(_05094_),
    .Y(_05095_)
  );
  sg13g2_o21ai_1 _15103_ (
    .A1(_00899_),
    .A2(_00651_),
    .B1(_01481_),
    .Y(_05096_)
  );
  sg13g2_a21oi_1 _15104_ (
    .A1(addr_i_7_),
    .A2(_02165_),
    .B1(_01514_),
    .Y(_05097_)
  );
  sg13g2_a21oi_1 _15105_ (
    .A1(addr_i_3_),
    .A2(_05096_),
    .B1(_05097_),
    .Y(_05098_)
  );
  sg13g2_o21ai_1 _15106_ (
    .A1(_00807_),
    .A2(_05098_),
    .B1(addr_i_11_),
    .Y(_05099_)
  );
  sg13g2_a21o_1 _15107_ (
    .A1(_05074_),
    .A2(_05095_),
    .B1(_05099_),
    .X(_05100_)
  );
  sg13g2_o21ai_1 _15108_ (
    .A1(_05000_),
    .A2(_05071_),
    .B1(_05100_),
    .Y(_05101_)
  );
  sg13g2_nor2_1 _15109_ (
    .A(_01526_),
    .B(_00923_),
    .Y(_05102_)
  );
  sg13g2_nor2_1 _15110_ (
    .A(_01616_),
    .B(_05102_),
    .Y(_05104_)
  );
  sg13g2_nand2_1 _15111_ (
    .A(_01917_),
    .B(_00607_),
    .Y(_05105_)
  );
  sg13g2_o21ai_1 _15112_ (
    .A1(addr_i_3_),
    .A2(_05104_),
    .B1(_05105_),
    .Y(_05106_)
  );
  sg13g2_nand2_1 _15113_ (
    .A(addr_i_5_),
    .B(_01933_),
    .Y(_05107_)
  );
  sg13g2_o21ai_1 _15114_ (
    .A1(addr_i_5_),
    .A2(_06021_),
    .B1(addr_i_3_),
    .Y(_05108_)
  );
  sg13g2_a21oi_1 _15115_ (
    .A1(_05107_),
    .A2(_05108_),
    .B1(addr_i_2_),
    .Y(_05109_)
  );
  sg13g2_a21oi_1 _15116_ (
    .A1(addr_i_2_),
    .A2(_05106_),
    .B1(_05109_),
    .Y(_05110_)
  );
  sg13g2_a22oi_1 _15117_ (
    .A1(addr_i_8_),
    .A2(_00184_),
    .B1(_01923_),
    .B2(_01169_),
    .Y(_05111_)
  );
  sg13g2_nor2b_1 _15118_ (
    .A(addr_i_8_),
    .B_N(addr_i_2_),
    .Y(_05112_)
  );
  sg13g2_nor3_1 _15119_ (
    .A(addr_i_3_),
    .B(_00128_),
    .C(_05112_),
    .Y(_05113_)
  );
  sg13g2_o21ai_1 _15120_ (
    .A1(_05111_),
    .A2(_05113_),
    .B1(_01937_),
    .Y(_05115_)
  );
  sg13g2_nand2_1 _15121_ (
    .A(addr_i_8_),
    .B(_04860_),
    .Y(_05116_)
  );
  sg13g2_a21oi_1 _15122_ (
    .A1(_02781_),
    .A2(_05116_),
    .B1(_00703_),
    .Y(_05117_)
  );
  sg13g2_a22oi_1 _15123_ (
    .A1(addr_i_4_),
    .A2(_05115_),
    .B1(_05117_),
    .B2(addr_i_7_),
    .Y(_05118_)
  );
  sg13g2_o21ai_1 _15124_ (
    .A1(addr_i_4_),
    .A2(_05110_),
    .B1(_05118_),
    .Y(_05119_)
  );
  sg13g2_a21oi_1 _15125_ (
    .A1(addr_i_2_),
    .A2(_01917_),
    .B1(_01031_),
    .Y(_05120_)
  );
  sg13g2_nor2_1 _15126_ (
    .A(_08410_),
    .B(_01911_),
    .Y(_05121_)
  );
  sg13g2_a21oi_1 _15127_ (
    .A1(_00170_),
    .A2(_01656_),
    .B1(_05121_),
    .Y(_05122_)
  );
  sg13g2_o21ai_1 _15128_ (
    .A1(addr_i_5_),
    .A2(_05120_),
    .B1(_05122_),
    .Y(_05123_)
  );
  sg13g2_a21oi_1 _15129_ (
    .A1(addr_i_6_),
    .A2(_03465_),
    .B1(addr_i_3_),
    .Y(_05124_)
  );
  sg13g2_o21ai_1 _15130_ (
    .A1(_05102_),
    .A2(_05124_),
    .B1(_01520_),
    .Y(_05126_)
  );
  sg13g2_nor2_1 _15131_ (
    .A(_03930_),
    .B(_02143_),
    .Y(_05127_)
  );
  sg13g2_a22oi_1 _15132_ (
    .A1(_00157_),
    .A2(_01923_),
    .B1(addr_i_2_),
    .B2(_06408_),
    .Y(_05128_)
  );
  sg13g2_a21oi_1 _15133_ (
    .A1(_05126_),
    .A2(_05127_),
    .B1(_05128_),
    .Y(_05129_)
  );
  sg13g2_a21oi_1 _15134_ (
    .A1(_01559_),
    .A2(_00500_),
    .B1(_03619_),
    .Y(_05130_)
  );
  sg13g2_o21ai_1 _15135_ (
    .A1(addr_i_5_),
    .A2(_05130_),
    .B1(addr_i_7_),
    .Y(_05131_)
  );
  sg13g2_a22oi_1 _15136_ (
    .A1(addr_i_3_),
    .A2(_05123_),
    .B1(_05129_),
    .B2(_05131_),
    .Y(_05132_)
  );
  sg13g2_nor2_1 _15137_ (
    .A(_01452_),
    .B(_05132_),
    .Y(_05133_)
  );
  sg13g2_a21oi_1 _15138_ (
    .A1(addr_i_6_),
    .A2(_02165_),
    .B1(addr_i_8_),
    .Y(_05134_)
  );
  sg13g2_o21ai_1 _15139_ (
    .A1(addr_i_2_),
    .A2(_06320_),
    .B1(_01570_),
    .Y(_05135_)
  );
  sg13g2_a21oi_1 _15140_ (
    .A1(addr_i_3_),
    .A2(_05135_),
    .B1(_06441_),
    .Y(_05137_)
  );
  sg13g2_a21oi_1 _15141_ (
    .A1(_00413_),
    .A2(_03465_),
    .B1(addr_i_3_),
    .Y(_05138_)
  );
  sg13g2_nand3b_1 _15142_ (
    .A_N(addr_i_5_),
    .B(addr_i_6_),
    .C(addr_i_8_),
    .Y(_05139_)
  );
  sg13g2_a21oi_1 _15143_ (
    .A1(_00915_),
    .A2(_05139_),
    .B1(_02343_),
    .Y(_05140_)
  );
  sg13g2_o21ai_1 _15144_ (
    .A1(_05138_),
    .A2(_05140_),
    .B1(addr_i_4_),
    .Y(_05141_)
  );
  sg13g2_o21ai_1 _15145_ (
    .A1(addr_i_4_),
    .A2(_05137_),
    .B1(_05141_),
    .Y(_05142_)
  );
  sg13g2_a22oi_1 _15146_ (
    .A1(_07824_),
    .A2(_06320_),
    .B1(_05134_),
    .B2(_05142_),
    .Y(_05143_)
  );
  sg13g2_nor3_1 _15147_ (
    .A(_01548_),
    .B(_00549_),
    .C(_00534_),
    .Y(_05144_)
  );
  sg13g2_o21ai_1 _15148_ (
    .A1(_05112_),
    .A2(_05144_),
    .B1(addr_i_3_),
    .Y(_05145_)
  );
  sg13g2_nor2_1 _15149_ (
    .A(_06198_),
    .B(_01252_),
    .Y(_05146_)
  );
  sg13g2_a21oi_1 _15150_ (
    .A1(_00549_),
    .A2(_01933_),
    .B1(addr_i_3_),
    .Y(_05148_)
  );
  sg13g2_o21ai_1 _15151_ (
    .A1(_05146_),
    .A2(_05148_),
    .B1(_03263_),
    .Y(_05149_)
  );
  sg13g2_nand3_1 _15152_ (
    .A(addr_i_5_),
    .B(_01933_),
    .C(_02781_),
    .Y(_05150_)
  );
  sg13g2_a21oi_1 _15153_ (
    .A1(_01729_),
    .A2(_05150_),
    .B1(_06419_),
    .Y(_05151_)
  );
  sg13g2_a22oi_1 _15154_ (
    .A1(_03465_),
    .A2(_02781_),
    .B1(addr_i_3_),
    .B2(addr_i_2_),
    .Y(_05152_)
  );
  sg13g2_o21ai_1 _15155_ (
    .A1(_05151_),
    .A2(_05152_),
    .B1(_00360_),
    .Y(_05153_)
  );
  sg13g2_a21oi_1 _15156_ (
    .A1(_00561_),
    .A2(_05112_),
    .B1(_06619_),
    .Y(_05154_)
  );
  sg13g2_nand4_1 _15157_ (
    .A(_05145_),
    .B(_05149_),
    .C(_05153_),
    .D(_05154_),
    .Y(_05155_)
  );
  sg13g2_o21ai_1 _15158_ (
    .A1(addr_i_7_),
    .A2(_05143_),
    .B1(_05155_),
    .Y(_05156_)
  );
  sg13g2_a21o_1 _15159_ (
    .A1(_00773_),
    .A2(_05156_),
    .B1(addr_i_11_),
    .X(_05157_)
  );
  sg13g2_a21oi_1 _15160_ (
    .A1(_00571_),
    .A2(_00878_),
    .B1(_00463_),
    .Y(_05159_)
  );
  sg13g2_a21oi_1 _15161_ (
    .A1(_02602_),
    .A2(_02887_),
    .B1(_00120_),
    .Y(_05160_)
  );
  sg13g2_or4_1 _15162_ (
    .A(_08332_),
    .B(_02361_),
    .C(_05159_),
    .D(_05160_),
    .X(_05161_)
  );
  sg13g2_a21oi_1 _15163_ (
    .A1(addr_i_6_),
    .A2(_01672_),
    .B1(_00844_),
    .Y(_05162_)
  );
  sg13g2_o21ai_1 _15164_ (
    .A1(_08410_),
    .A2(_05162_),
    .B1(addr_i_3_),
    .Y(_05163_)
  );
  sg13g2_a21oi_1 _15165_ (
    .A1(_00065_),
    .A2(_00819_),
    .B1(_00648_),
    .Y(_05164_)
  );
  sg13g2_o21ai_1 _15166_ (
    .A1(_01064_),
    .A2(_05164_),
    .B1(_04251_),
    .Y(_05165_)
  );
  sg13g2_nand4_1 _15167_ (
    .A(_00629_),
    .B(_05161_),
    .C(_05163_),
    .D(_05165_),
    .Y(_05166_)
  );
  sg13g2_nor2_1 _15168_ (
    .A(_08332_),
    .B(_01112_),
    .Y(_05167_)
  );
  sg13g2_a221oi_1 _15169_ (
    .A1(addr_i_4_),
    .A2(_00473_),
    .B1(_01254_),
    .B2(addr_i_5_),
    .C1(addr_i_7_),
    .Y(_05168_)
  );
  sg13g2_a22oi_1 _15170_ (
    .A1(_00815_),
    .A2(_05167_),
    .B1(_05168_),
    .B2(_00485_),
    .Y(_05171_)
  );
  sg13g2_o21ai_1 _15171_ (
    .A1(addr_i_6_),
    .A2(_06220_),
    .B1(_03809_),
    .Y(_05172_)
  );
  sg13g2_a21oi_1 _15172_ (
    .A1(_00032_),
    .A2(_05172_),
    .B1(_08000_),
    .Y(_05173_)
  );
  sg13g2_o21ai_1 _15173_ (
    .A1(_00654_),
    .A2(_05173_),
    .B1(_00565_),
    .Y(_05174_)
  );
  sg13g2_a21oi_1 _15174_ (
    .A1(_09415_),
    .A2(_00037_),
    .B1(addr_i_4_),
    .Y(_05175_)
  );
  sg13g2_a22oi_1 _15175_ (
    .A1(_02268_),
    .A2(_01228_),
    .B1(_05175_),
    .B2(_05888_),
    .Y(_05176_)
  );
  sg13g2_nand3b_1 _15176_ (
    .A_N(_05171_),
    .B(_05174_),
    .C(_05176_),
    .Y(_05177_)
  );
  sg13g2_and2_1 _15177_ (
    .A(_05166_),
    .B(_05177_),
    .X(_05178_)
  );
  sg13g2_nor3_1 _15178_ (
    .A(_03455_),
    .B(_00667_),
    .C(_02226_),
    .Y(_05179_)
  );
  sg13g2_a21oi_1 _15179_ (
    .A1(addr_i_5_),
    .A2(_05910_),
    .B1(addr_i_3_),
    .Y(_05180_)
  );
  sg13g2_o21ai_1 _15180_ (
    .A1(_07879_),
    .A2(_05180_),
    .B1(addr_i_2_),
    .Y(_05182_)
  );
  sg13g2_a21oi_1 _15181_ (
    .A1(_00238_),
    .A2(_00786_),
    .B1(_03632_),
    .Y(_05183_)
  );
  sg13g2_a21oi_1 _15182_ (
    .A1(_05182_),
    .A2(_05183_),
    .B1(addr_i_7_),
    .Y(_05184_)
  );
  sg13g2_a21oi_1 _15183_ (
    .A1(_07569_),
    .A2(_01894_),
    .B1(_02759_),
    .Y(_05185_)
  );
  sg13g2_a22oi_1 _15184_ (
    .A1(_01320_),
    .A2(_05179_),
    .B1(_05184_),
    .B2(_05185_),
    .Y(_05186_)
  );
  sg13g2_nand2_1 _15185_ (
    .A(_01008_),
    .B(_04881_),
    .Y(_05187_)
  );
  sg13g2_o21ai_1 _15186_ (
    .A1(_01200_),
    .A2(_05187_),
    .B1(addr_i_5_),
    .Y(_05188_)
  );
  sg13g2_o21ai_1 _15187_ (
    .A1(_01659_),
    .A2(_02441_),
    .B1(addr_i_3_),
    .Y(_05189_)
  );
  sg13g2_o21ai_1 _15188_ (
    .A1(_05037_),
    .A2(_04490_),
    .B1(addr_i_6_),
    .Y(_05190_)
  );
  sg13g2_a21oi_1 _15189_ (
    .A1(_05189_),
    .A2(_05190_),
    .B1(_06619_),
    .Y(_05191_)
  );
  sg13g2_a21oi_1 _15190_ (
    .A1(_01008_),
    .A2(_00405_),
    .B1(_00697_),
    .Y(_05193_)
  );
  sg13g2_o21ai_1 _15191_ (
    .A1(_00090_),
    .A2(_03570_),
    .B1(addr_i_8_),
    .Y(_05194_)
  );
  sg13g2_nor2_1 _15192_ (
    .A(_04075_),
    .B(_08941_),
    .Y(_05195_)
  );
  sg13g2_nor4_1 _15193_ (
    .A(_01155_),
    .B(_08598_),
    .C(_00009_),
    .D(_05195_),
    .Y(_05196_)
  );
  sg13g2_nor4_1 _15194_ (
    .A(_05191_),
    .B(_05193_),
    .C(_05194_),
    .D(_05196_),
    .Y(_05197_)
  );
  sg13g2_a221oi_1 _15195_ (
    .A1(_01151_),
    .A2(_05186_),
    .B1(_05188_),
    .B2(_05197_),
    .C1(addr_i_9_),
    .Y(_05198_)
  );
  sg13g2_a22oi_1 _15196_ (
    .A1(addr_i_9_),
    .A2(_05178_),
    .B1(_05198_),
    .B2(_00511_),
    .Y(_05199_)
  );
  sg13g2_a22oi_1 _15197_ (
    .A1(_05119_),
    .A2(_05133_),
    .B1(_05157_),
    .B2(_05199_),
    .Y(_05200_)
  );
  sg13g2_a21oi_1 _15198_ (
    .A1(_02528_),
    .A2(_01704_),
    .B1(_00701_),
    .Y(_05201_)
  );
  sg13g2_a22oi_1 _15199_ (
    .A1(_00073_),
    .A2(_03723_),
    .B1(_05201_),
    .B2(_01324_),
    .Y(_05202_)
  );
  sg13g2_a21oi_1 _15200_ (
    .A1(_00476_),
    .A2(_00376_),
    .B1(addr_i_3_),
    .Y(_05204_)
  );
  sg13g2_o21ai_1 _15201_ (
    .A1(addr_i_4_),
    .A2(_01326_),
    .B1(_05204_),
    .Y(_05205_)
  );
  sg13g2_o21ai_1 _15202_ (
    .A1(_00010_),
    .A2(_00384_),
    .B1(_03281_),
    .Y(_05206_)
  );
  sg13g2_nand3_1 _15203_ (
    .A(addr_i_3_),
    .B(_04087_),
    .C(_05206_),
    .Y(_05207_)
  );
  sg13g2_a21oi_1 _15204_ (
    .A1(_05205_),
    .A2(_05207_),
    .B1(addr_i_5_),
    .Y(_05208_)
  );
  sg13g2_a21oi_1 _15205_ (
    .A1(_07204_),
    .A2(_00878_),
    .B1(_05822_),
    .Y(_05209_)
  );
  sg13g2_a22oi_1 _15206_ (
    .A1(_01508_),
    .A2(_04786_),
    .B1(_05209_),
    .B2(addr_i_8_),
    .Y(_05210_)
  );
  sg13g2_o21ai_1 _15207_ (
    .A1(_05202_),
    .A2(_05208_),
    .B1(_05210_),
    .Y(_05211_)
  );
  sg13g2_o21ai_1 _15208_ (
    .A1(addr_i_7_),
    .A2(_01276_),
    .B1(_08166_),
    .Y(_05212_)
  );
  sg13g2_o21ai_1 _15209_ (
    .A1(_00914_),
    .A2(_01572_),
    .B1(_05212_),
    .Y(_05213_)
  );
  sg13g2_o21ai_1 _15210_ (
    .A1(_03577_),
    .A2(_05213_),
    .B1(addr_i_3_),
    .Y(_05215_)
  );
  sg13g2_nor3_1 _15211_ (
    .A(addr_i_6_),
    .B(_00269_),
    .C(_00400_),
    .Y(_05216_)
  );
  sg13g2_a21oi_1 _15212_ (
    .A1(_01077_),
    .A2(_05689_),
    .B1(addr_i_3_),
    .Y(_05217_)
  );
  sg13g2_buf_1 _15213_ (
    .A(_03809_),
    .X(_05218_)
  );
  sg13g2_o21ai_1 _15214_ (
    .A1(_05216_),
    .A2(_05217_),
    .B1(_05218_),
    .Y(_05219_)
  );
  sg13g2_nor2_1 _15215_ (
    .A(_03776_),
    .B(_03245_),
    .Y(_05220_)
  );
  sg13g2_o21ai_1 _15216_ (
    .A1(_00384_),
    .A2(_00031_),
    .B1(_05220_),
    .Y(_05221_)
  );
  sg13g2_nand4_1 _15217_ (
    .A(addr_i_8_),
    .B(_05215_),
    .C(_05219_),
    .D(_05221_),
    .Y(_05222_)
  );
  sg13g2_and2_1 _15218_ (
    .A(addr_i_10_),
    .B(_05222_),
    .X(_05223_)
  );
  sg13g2_a21oi_1 _15219_ (
    .A1(_05211_),
    .A2(_05223_),
    .B1(addr_i_9_),
    .Y(_05224_)
  );
  sg13g2_nand2b_1 _15220_ (
    .A_N(_00023_),
    .B(_01234_),
    .Y(_05226_)
  );
  sg13g2_a21oi_1 _15221_ (
    .A1(_02815_),
    .A2(_01622_),
    .B1(_02191_),
    .Y(_05227_)
  );
  sg13g2_a21oi_1 _15222_ (
    .A1(_00838_),
    .A2(_01990_),
    .B1(_05227_),
    .Y(_05228_)
  );
  sg13g2_a21oi_1 _15223_ (
    .A1(_00056_),
    .A2(_05228_),
    .B1(addr_i_3_),
    .Y(_05229_)
  );
  sg13g2_o21ai_1 _15224_ (
    .A1(addr_i_7_),
    .A2(_03150_),
    .B1(addr_i_3_),
    .Y(_05230_)
  );
  sg13g2_nor2_1 _15225_ (
    .A(addr_i_5_),
    .B(_05225_),
    .Y(_05231_)
  );
  sg13g2_nor2_1 _15226_ (
    .A(_02577_),
    .B(_00522_),
    .Y(_05232_)
  );
  sg13g2_a21oi_1 _15227_ (
    .A1(addr_i_4_),
    .A2(_05231_),
    .B1(_05232_),
    .Y(_05233_)
  );
  sg13g2_a21oi_1 _15228_ (
    .A1(_05230_),
    .A2(_05233_),
    .B1(_00123_),
    .Y(_05234_)
  );
  sg13g2_a22oi_1 _15229_ (
    .A1(addr_i_4_),
    .A2(_05226_),
    .B1(_05229_),
    .B2(_05234_),
    .Y(_05235_)
  );
  sg13g2_nand2_1 _15230_ (
    .A(addr_i_4_),
    .B(_00435_),
    .Y(_05237_)
  );
  sg13g2_nand2_1 _15231_ (
    .A(addr_i_4_),
    .B(_01054_),
    .Y(_05238_)
  );
  sg13g2_a21oi_1 _15232_ (
    .A1(_00249_),
    .A2(_05238_),
    .B1(addr_i_6_),
    .Y(_05239_)
  );
  sg13g2_a21oi_1 _15233_ (
    .A1(_01104_),
    .A2(_02294_),
    .B1(addr_i_4_),
    .Y(_05240_)
  );
  sg13g2_a22oi_1 _15234_ (
    .A1(_00015_),
    .A2(_05237_),
    .B1(_05239_),
    .B2(_05240_),
    .Y(_05241_)
  );
  sg13g2_nand3_1 _15235_ (
    .A(_00122_),
    .B(_03325_),
    .C(_04077_),
    .Y(_05242_)
  );
  sg13g2_nor2_1 _15236_ (
    .A(_00120_),
    .B(_06220_),
    .Y(_05243_)
  );
  sg13g2_a21oi_1 _15237_ (
    .A1(_03226_),
    .A2(_05243_),
    .B1(_04068_),
    .Y(_05244_)
  );
  sg13g2_a21oi_1 _15238_ (
    .A1(_01301_),
    .A2(_01589_),
    .B1(addr_i_7_),
    .Y(_05245_)
  );
  sg13g2_a22oi_1 _15239_ (
    .A1(_05242_),
    .A2(_05244_),
    .B1(_05245_),
    .B2(addr_i_3_),
    .Y(_05246_)
  );
  sg13g2_a22oi_1 _15240_ (
    .A1(addr_i_3_),
    .A2(_05241_),
    .B1(_05246_),
    .B2(_07293_),
    .Y(_05248_)
  );
  sg13g2_nor2_1 _15241_ (
    .A(addr_i_10_),
    .B(_05248_),
    .Y(_05249_)
  );
  sg13g2_o21ai_1 _15242_ (
    .A1(addr_i_8_),
    .A2(_05235_),
    .B1(_05249_),
    .Y(_05250_)
  );
  sg13g2_o21ai_1 _15243_ (
    .A1(_05546_),
    .A2(_05231_),
    .B1(_01692_),
    .Y(_05251_)
  );
  sg13g2_nor2_1 _15244_ (
    .A(addr_i_4_),
    .B(_07038_),
    .Y(_05252_)
  );
  sg13g2_o21ai_1 _15245_ (
    .A1(_01402_),
    .A2(_05252_),
    .B1(addr_i_2_),
    .Y(_05253_)
  );
  sg13g2_nand2b_1 _15246_ (
    .A_N(_05251_),
    .B(_05253_),
    .Y(_05254_)
  );
  sg13g2_nand2_1 _15247_ (
    .A(_00010_),
    .B(_02107_),
    .Y(_05255_)
  );
  sg13g2_nand4_1 _15248_ (
    .A(_01199_),
    .B(_01704_),
    .C(_00852_),
    .D(_05255_),
    .Y(_05256_)
  );
  sg13g2_nand2_1 _15249_ (
    .A(_09459_),
    .B(_00783_),
    .Y(_05257_)
  );
  sg13g2_o21ai_1 _15250_ (
    .A1(_00959_),
    .A2(_09459_),
    .B1(_00375_),
    .Y(_05259_)
  );
  sg13g2_nand3_1 _15251_ (
    .A(_05257_),
    .B(_02315_),
    .C(_05259_),
    .Y(_05260_)
  );
  sg13g2_a221oi_1 _15252_ (
    .A1(_03260_),
    .A2(_05254_),
    .B1(_05256_),
    .B2(addr_i_5_),
    .C1(_05260_),
    .Y(_05261_)
  );
  sg13g2_o21ai_1 _15253_ (
    .A1(_08410_),
    .A2(_02042_),
    .B1(addr_i_3_),
    .Y(_05262_)
  );
  sg13g2_o21ai_1 _15254_ (
    .A1(addr_i_5_),
    .A2(_05943_),
    .B1(addr_i_4_),
    .Y(_05263_)
  );
  sg13g2_nand4_1 _15255_ (
    .A(_01118_),
    .B(_01524_),
    .C(_05262_),
    .D(_05263_),
    .Y(_05264_)
  );
  sg13g2_a221oi_1 _15256_ (
    .A1(_01292_),
    .A2(_08111_),
    .B1(_01439_),
    .B2(_01472_),
    .C1(_01049_),
    .Y(_05265_)
  );
  sg13g2_nor2_1 _15257_ (
    .A(_00030_),
    .B(_01406_),
    .Y(_05266_)
  );
  sg13g2_nor2_1 _15258_ (
    .A(_08299_),
    .B(_05266_),
    .Y(_05267_)
  );
  sg13g2_a21o_1 _15259_ (
    .A1(_05265_),
    .A2(_05267_),
    .B1(_07514_),
    .X(_05268_)
  );
  sg13g2_and2_1 _15260_ (
    .A(_05264_),
    .B(_05268_),
    .X(_05270_)
  );
  sg13g2_o21ai_1 _15261_ (
    .A1(addr_i_8_),
    .A2(_05261_),
    .B1(_05270_),
    .Y(_05271_)
  );
  sg13g2_o21ai_1 _15262_ (
    .A1(addr_i_2_),
    .A2(_01718_),
    .B1(_01065_),
    .Y(_05272_)
  );
  sg13g2_a21oi_1 _15263_ (
    .A1(_00695_),
    .A2(_01967_),
    .B1(_03281_),
    .Y(_05273_)
  );
  sg13g2_a21oi_1 _15264_ (
    .A1(addr_i_4_),
    .A2(_05272_),
    .B1(_05273_),
    .Y(_05274_)
  );
  sg13g2_a221oi_1 _15265_ (
    .A1(_05745_),
    .A2(_06298_),
    .B1(_00442_),
    .B2(_04092_),
    .C1(addr_i_7_),
    .Y(_05275_)
  );
  sg13g2_a22oi_1 _15266_ (
    .A1(_00120_),
    .A2(_00550_),
    .B1(_06563_),
    .B2(addr_i_4_),
    .Y(_05276_)
  );
  sg13g2_a221oi_1 _15267_ (
    .A1(_00260_),
    .A2(_00676_),
    .B1(_05379_),
    .B2(_07326_),
    .C1(_00956_),
    .Y(_05277_)
  );
  sg13g2_o21ai_1 _15268_ (
    .A1(_05276_),
    .A2(_05277_),
    .B1(addr_i_7_),
    .Y(_05278_)
  );
  sg13g2_nand2b_1 _15269_ (
    .A_N(_05275_),
    .B(_05278_),
    .Y(_05279_)
  );
  sg13g2_o21ai_1 _15270_ (
    .A1(addr_i_3_),
    .A2(_05274_),
    .B1(_05279_),
    .Y(_05282_)
  );
  sg13g2_a21oi_1 _15271_ (
    .A1(_03347_),
    .A2(_00037_),
    .B1(addr_i_4_),
    .Y(_05283_)
  );
  sg13g2_o21ai_1 _15272_ (
    .A1(_04915_),
    .A2(_05283_),
    .B1(_00949_),
    .Y(_05284_)
  );
  sg13g2_and2_1 _15273_ (
    .A(_06695_),
    .B(_05284_),
    .X(_05285_)
  );
  sg13g2_o21ai_1 _15274_ (
    .A1(_00322_),
    .A2(_01450_),
    .B1(addr_i_4_),
    .Y(_05286_)
  );
  sg13g2_o21ai_1 _15275_ (
    .A1(addr_i_3_),
    .A2(_03485_),
    .B1(_05286_),
    .Y(_05287_)
  );
  sg13g2_a21oi_1 _15276_ (
    .A1(addr_i_3_),
    .A2(_02119_),
    .B1(_00990_),
    .Y(_05288_)
  );
  sg13g2_nor2_1 _15277_ (
    .A(addr_i_7_),
    .B(_05288_),
    .Y(_05289_)
  );
  sg13g2_a21oi_1 _15278_ (
    .A1(_00981_),
    .A2(_04093_),
    .B1(_02803_),
    .Y(_05290_)
  );
  sg13g2_a22oi_1 _15279_ (
    .A1(addr_i_7_),
    .A2(_05287_),
    .B1(_05289_),
    .B2(_05290_),
    .Y(_05291_)
  );
  sg13g2_a221oi_1 _15280_ (
    .A1(addr_i_8_),
    .A2(_05282_),
    .B1(_05285_),
    .B2(_05291_),
    .C1(addr_i_10_),
    .Y(_05293_)
  );
  sg13g2_a22oi_1 _15281_ (
    .A1(addr_i_10_),
    .A2(_05271_),
    .B1(_05293_),
    .B2(_00397_),
    .Y(_05294_)
  );
  sg13g2_a22oi_1 _15282_ (
    .A1(_05224_),
    .A2(_05250_),
    .B1(_01640_),
    .B2(_05294_),
    .Y(_05295_)
  );
  sg13g2_o21ai_1 _15283_ (
    .A1(_05200_),
    .A2(_05295_),
    .B1(_02251_),
    .Y(_05296_)
  );
  sg13g2_o21ai_1 _15284_ (
    .A1(_02251_),
    .A2(_05101_),
    .B1(_05296_),
    .Y(data_o_23_)
  );
  sg13g2_a21oi_1 _15285_ (
    .A1(addr_i_3_),
    .A2(_01493_),
    .B1(_02265_),
    .Y(_05297_)
  );
  sg13g2_nor2_1 _15286_ (
    .A(_03292_),
    .B(_07348_),
    .Y(_05298_)
  );
  sg13g2_nor2_1 _15287_ (
    .A(_07237_),
    .B(_03106_),
    .Y(_05299_)
  );
  sg13g2_nor2_1 _15288_ (
    .A(_02086_),
    .B(_05299_),
    .Y(_05300_)
  );
  sg13g2_nor3_1 _15289_ (
    .A(addr_i_2_),
    .B(_00009_),
    .C(_05300_),
    .Y(_05301_)
  );
  sg13g2_a22oi_1 _15290_ (
    .A1(_05297_),
    .A2(_05298_),
    .B1(_05301_),
    .B2(_03494_),
    .Y(_05303_)
  );
  sg13g2_nand2_1 _15291_ (
    .A(addr_i_5_),
    .B(_08774_),
    .Y(_05304_)
  );
  sg13g2_o21ai_1 _15292_ (
    .A1(addr_i_3_),
    .A2(_05304_),
    .B1(_00328_),
    .Y(_05305_)
  );
  sg13g2_nor2_1 _15293_ (
    .A(addr_i_4_),
    .B(_02672_),
    .Y(_05306_)
  );
  sg13g2_a221oi_1 _15294_ (
    .A1(addr_i_3_),
    .A2(_05304_),
    .B1(_05305_),
    .B2(addr_i_4_),
    .C1(_05306_),
    .Y(_05307_)
  );
  sg13g2_nor2_1 _15295_ (
    .A(_02535_),
    .B(_05307_),
    .Y(_05308_)
  );
  sg13g2_o21ai_1 _15296_ (
    .A1(addr_i_2_),
    .A2(_01439_),
    .B1(_08232_),
    .Y(_05309_)
  );
  sg13g2_a21oi_1 _15297_ (
    .A1(_03540_),
    .A2(_01658_),
    .B1(_08951_),
    .Y(_05310_)
  );
  sg13g2_a21o_1 _15298_ (
    .A1(_01131_),
    .A2(_05309_),
    .B1(_05310_),
    .X(_05311_)
  );
  sg13g2_a21oi_1 _15299_ (
    .A1(_01967_),
    .A2(_03346_),
    .B1(addr_i_5_),
    .Y(_05312_)
  );
  sg13g2_a21oi_1 _15300_ (
    .A1(_03424_),
    .A2(_00317_),
    .B1(addr_i_3_),
    .Y(_05314_)
  );
  sg13g2_a22oi_1 _15301_ (
    .A1(addr_i_5_),
    .A2(_05311_),
    .B1(_05312_),
    .B2(_05314_),
    .Y(_05315_)
  );
  sg13g2_o21ai_1 _15302_ (
    .A1(_01612_),
    .A2(_05315_),
    .B1(_01773_),
    .Y(_05316_)
  );
  sg13g2_nor3_1 _15303_ (
    .A(_05303_),
    .B(_05308_),
    .C(_05316_),
    .Y(_05317_)
  );
  sg13g2_o21ai_1 _15304_ (
    .A1(_00742_),
    .A2(_00890_),
    .B1(addr_i_4_),
    .Y(_05318_)
  );
  sg13g2_a21oi_1 _15305_ (
    .A1(_02497_),
    .A2(_05318_),
    .B1(addr_i_7_),
    .Y(_05319_)
  );
  sg13g2_nand3_1 _15306_ (
    .A(_02777_),
    .B(_01065_),
    .C(_00244_),
    .Y(_05320_)
  );
  sg13g2_nand2_1 _15307_ (
    .A(_04741_),
    .B(_05320_),
    .Y(_05321_)
  );
  sg13g2_o21ai_1 _15308_ (
    .A1(_05319_),
    .A2(_05321_),
    .B1(_03260_),
    .Y(_05322_)
  );
  sg13g2_a21o_1 _15309_ (
    .A1(addr_i_2_),
    .A2(_01154_),
    .B1(_08299_),
    .X(_05323_)
  );
  sg13g2_o21ai_1 _15310_ (
    .A1(addr_i_7_),
    .A2(_09497_),
    .B1(_00065_),
    .Y(_05325_)
  );
  sg13g2_a22oi_1 _15311_ (
    .A1(_00871_),
    .A2(_05325_),
    .B1(_00799_),
    .B2(addr_i_6_),
    .Y(_05326_)
  );
  sg13g2_a221oi_1 _15312_ (
    .A1(_02277_),
    .A2(_04982_),
    .B1(_05323_),
    .B2(_00258_),
    .C1(_05326_),
    .Y(_05327_)
  );
  sg13g2_a21o_1 _15313_ (
    .A1(_05322_),
    .A2(_05327_),
    .B1(_07293_),
    .X(_05328_)
  );
  sg13g2_nor3_1 _15314_ (
    .A(addr_i_6_),
    .B(_01019_),
    .C(_07337_),
    .Y(_05329_)
  );
  sg13g2_nand2_1 _15315_ (
    .A(_00115_),
    .B(_02785_),
    .Y(_05330_)
  );
  sg13g2_a21oi_1 _15316_ (
    .A1(_04379_),
    .A2(_05330_),
    .B1(addr_i_5_),
    .Y(_05331_)
  );
  sg13g2_o21ai_1 _15317_ (
    .A1(_05329_),
    .A2(_05331_),
    .B1(_00779_),
    .Y(_05332_)
  );
  sg13g2_nand2_1 _15318_ (
    .A(addr_i_2_),
    .B(_01636_),
    .Y(_05333_)
  );
  sg13g2_nand2_1 _15319_ (
    .A(addr_i_3_),
    .B(_05333_),
    .Y(_05334_)
  );
  sg13g2_nand4_1 _15320_ (
    .A(_07337_),
    .B(_09138_),
    .C(_00545_),
    .D(_05334_),
    .Y(_05336_)
  );
  sg13g2_nor3_1 _15321_ (
    .A(_00548_),
    .B(_02241_),
    .C(_04261_),
    .Y(_05337_)
  );
  sg13g2_a22oi_1 _15322_ (
    .A1(_01355_),
    .A2(_04499_),
    .B1(_05337_),
    .B2(addr_i_8_),
    .Y(_05338_)
  );
  sg13g2_nand3_1 _15323_ (
    .A(_05332_),
    .B(_05336_),
    .C(_05338_),
    .Y(_05339_)
  );
  sg13g2_nand3_1 _15324_ (
    .A(addr_i_9_),
    .B(_05328_),
    .C(_05339_),
    .Y(_05340_)
  );
  sg13g2_o21ai_1 _15325_ (
    .A1(_07248_),
    .A2(_08188_),
    .B1(addr_i_3_),
    .Y(_05341_)
  );
  sg13g2_o21ai_1 _15326_ (
    .A1(addr_i_7_),
    .A2(_00514_),
    .B1(_05341_),
    .Y(_05342_)
  );
  sg13g2_a21oi_1 _15327_ (
    .A1(_03292_),
    .A2(_05342_),
    .B1(_00081_),
    .Y(_05343_)
  );
  sg13g2_a21oi_1 _15328_ (
    .A1(addr_i_4_),
    .A2(_02135_),
    .B1(_01232_),
    .Y(_05344_)
  );
  sg13g2_nand2_1 _15329_ (
    .A(_01203_),
    .B(_01056_),
    .Y(_05345_)
  );
  sg13g2_a221oi_1 _15330_ (
    .A1(_01585_),
    .A2(_02304_),
    .B1(_05345_),
    .B2(addr_i_6_),
    .C1(addr_i_3_),
    .Y(_05347_)
  );
  sg13g2_a21o_1 _15331_ (
    .A1(addr_i_3_),
    .A2(_05344_),
    .B1(_05347_),
    .X(_05348_)
  );
  sg13g2_a21oi_1 _15332_ (
    .A1(_05343_),
    .A2(_05348_),
    .B1(_02368_),
    .Y(_05349_)
  );
  sg13g2_a21oi_1 _15333_ (
    .A1(_00820_),
    .A2(_00470_),
    .B1(_00409_),
    .Y(_05350_)
  );
  sg13g2_a22oi_1 _15334_ (
    .A1(_00115_),
    .A2(_03325_),
    .B1(_03348_),
    .B2(_03150_),
    .Y(_05351_)
  );
  sg13g2_nor2_1 _15335_ (
    .A(addr_i_2_),
    .B(_05351_),
    .Y(_05352_)
  );
  sg13g2_a22oi_1 _15336_ (
    .A1(addr_i_3_),
    .A2(_02342_),
    .B1(_05350_),
    .B2(_05352_),
    .Y(_05353_)
  );
  sg13g2_o21ai_1 _15337_ (
    .A1(_00022_),
    .A2(_03455_),
    .B1(addr_i_3_),
    .Y(_05354_)
  );
  sg13g2_o21ai_1 _15338_ (
    .A1(_08575_),
    .A2(_01845_),
    .B1(_02796_),
    .Y(_05355_)
  );
  sg13g2_nand4_1 _15339_ (
    .A(_01168_),
    .B(_03890_),
    .C(_05354_),
    .D(_05355_),
    .Y(_05356_)
  );
  sg13g2_o21ai_1 _15340_ (
    .A1(_02963_),
    .A2(_05353_),
    .B1(_05356_),
    .Y(_05358_)
  );
  sg13g2_a21oi_1 _15341_ (
    .A1(_00020_),
    .A2(_02076_),
    .B1(addr_i_4_),
    .Y(_05359_)
  );
  sg13g2_nor2_1 _15342_ (
    .A(_00007_),
    .B(_05359_),
    .Y(_05360_)
  );
  sg13g2_nor2_1 _15343_ (
    .A(addr_i_3_),
    .B(_04086_),
    .Y(_05361_)
  );
  sg13g2_xnor2_1 _15344_ (
    .A(addr_i_4_),
    .B(_05361_),
    .Y(_05362_)
  );
  sg13g2_a221oi_1 _15345_ (
    .A1(_09039_),
    .A2(_05360_),
    .B1(_05362_),
    .B2(_01320_),
    .C1(addr_i_8_),
    .Y(_05363_)
  );
  sg13g2_a21oi_1 _15346_ (
    .A1(addr_i_3_),
    .A2(_01301_),
    .B1(_07889_),
    .Y(_05364_)
  );
  sg13g2_nand2_1 _15347_ (
    .A(_00151_),
    .B(_01749_),
    .Y(_05365_)
  );
  sg13g2_a22oi_1 _15348_ (
    .A1(addr_i_5_),
    .A2(_05365_),
    .B1(_05932_),
    .B2(addr_i_7_),
    .Y(_05366_)
  );
  sg13g2_o21ai_1 _15349_ (
    .A1(addr_i_2_),
    .A2(_05364_),
    .B1(_05366_),
    .Y(_05367_)
  );
  sg13g2_o21ai_1 _15350_ (
    .A1(_01086_),
    .A2(_00177_),
    .B1(addr_i_3_),
    .Y(_05369_)
  );
  sg13g2_nand4_1 _15351_ (
    .A(_00138_),
    .B(_02047_),
    .C(_03827_),
    .D(_05369_),
    .Y(_05370_)
  );
  sg13g2_a22oi_1 _15352_ (
    .A1(addr_i_3_),
    .A2(_05333_),
    .B1(_00503_),
    .B2(_00268_),
    .Y(_05371_)
  );
  sg13g2_o21ai_1 _15353_ (
    .A1(_00317_),
    .A2(_05371_),
    .B1(addr_i_8_),
    .Y(_05372_)
  );
  sg13g2_nor2_1 _15354_ (
    .A(_00910_),
    .B(_04579_),
    .Y(_05373_)
  );
  sg13g2_nor3_1 _15355_ (
    .A(_00324_),
    .B(_01540_),
    .C(_05373_),
    .Y(_05374_)
  );
  sg13g2_a22oi_1 _15356_ (
    .A1(addr_i_7_),
    .A2(_05370_),
    .B1(_05372_),
    .B2(_05374_),
    .Y(_05375_)
  );
  sg13g2_a22oi_1 _15357_ (
    .A1(_05363_),
    .A2(_05367_),
    .B1(_00396_),
    .B2(_05375_),
    .Y(_05376_)
  );
  sg13g2_nor4_1 _15358_ (
    .A(_03841_),
    .B(_05349_),
    .C(_05358_),
    .D(_05376_),
    .Y(_05377_)
  );
  sg13g2_a21oi_1 _15359_ (
    .A1(_05317_),
    .A2(_05340_),
    .B1(_05377_),
    .Y(_05378_)
  );
  sg13g2_o21ai_1 _15360_ (
    .A1(_02268_),
    .A2(_06574_),
    .B1(_03263_),
    .Y(_05380_)
  );
  sg13g2_a21oi_1 _15361_ (
    .A1(_03527_),
    .A2(_05380_),
    .B1(addr_i_7_),
    .Y(_05381_)
  );
  sg13g2_o21ai_1 _15362_ (
    .A1(_00223_),
    .A2(_01481_),
    .B1(addr_i_4_),
    .Y(_05382_)
  );
  sg13g2_nand2b_1 _15363_ (
    .A_N(_05381_),
    .B(_05382_),
    .Y(_05383_)
  );
  sg13g2_nor2_1 _15364_ (
    .A(_00243_),
    .B(_02397_),
    .Y(_05384_)
  );
  sg13g2_o21ai_1 _15365_ (
    .A1(_09205_),
    .A2(_01901_),
    .B1(_07790_),
    .Y(_05385_)
  );
  sg13g2_nor2_1 _15366_ (
    .A(addr_i_5_),
    .B(_00968_),
    .Y(_05386_)
  );
  sg13g2_nor2_1 _15367_ (
    .A(_00261_),
    .B(_01421_),
    .Y(_05387_)
  );
  sg13g2_o21ai_1 _15368_ (
    .A1(_05386_),
    .A2(_05387_),
    .B1(addr_i_3_),
    .Y(_05388_)
  );
  sg13g2_o21ai_1 _15369_ (
    .A1(_01320_),
    .A2(_03433_),
    .B1(addr_i_2_),
    .Y(_05389_)
  );
  sg13g2_nand2_1 _15370_ (
    .A(_05388_),
    .B(_05389_),
    .Y(_05392_)
  );
  sg13g2_o21ai_1 _15371_ (
    .A1(_01616_),
    .A2(_00945_),
    .B1(_01240_),
    .Y(_05393_)
  );
  sg13g2_nand2_1 _15372_ (
    .A(_00423_),
    .B(_05393_),
    .Y(_05394_)
  );
  sg13g2_a221oi_1 _15373_ (
    .A1(addr_i_7_),
    .A2(_05385_),
    .B1(_05392_),
    .B2(addr_i_4_),
    .C1(_05394_),
    .Y(_05395_)
  );
  sg13g2_a22oi_1 _15374_ (
    .A1(_02604_),
    .A2(_05383_),
    .B1(_05384_),
    .B2(_05395_),
    .Y(_05396_)
  );
  sg13g2_a21oi_1 _15375_ (
    .A1(_06519_),
    .A2(_03084_),
    .B1(_03040_),
    .Y(_05397_)
  );
  sg13g2_o21ai_1 _15376_ (
    .A1(addr_i_10_),
    .A2(_05396_),
    .B1(_05397_),
    .Y(_05398_)
  );
  sg13g2_o21ai_1 _15377_ (
    .A1(addr_i_11_),
    .A2(_05378_),
    .B1(_05398_),
    .Y(_05399_)
  );
  sg13g2_o21ai_1 _15378_ (
    .A1(_00377_),
    .A2(_00617_),
    .B1(_01519_),
    .Y(_05400_)
  );
  sg13g2_nand2_1 _15379_ (
    .A(_04236_),
    .B(_05400_),
    .Y(_05401_)
  );
  sg13g2_a21oi_1 _15380_ (
    .A1(_00861_),
    .A2(_09507_),
    .B1(_06574_),
    .Y(_05403_)
  );
  sg13g2_o21ai_1 _15381_ (
    .A1(addr_i_4_),
    .A2(_05403_),
    .B1(_02406_),
    .Y(_05404_)
  );
  sg13g2_a21oi_1 _15382_ (
    .A1(_00927_),
    .A2(_09149_),
    .B1(_02777_),
    .Y(_05405_)
  );
  sg13g2_nand2_1 _15383_ (
    .A(addr_i_2_),
    .B(_05405_),
    .Y(_05406_)
  );
  sg13g2_o21ai_1 _15384_ (
    .A1(_00209_),
    .A2(_00301_),
    .B1(addr_i_3_),
    .Y(_05407_)
  );
  sg13g2_a21oi_1 _15385_ (
    .A1(_05406_),
    .A2(_05407_),
    .B1(_01095_),
    .Y(_05408_)
  );
  sg13g2_a22oi_1 _15386_ (
    .A1(_00123_),
    .A2(_05401_),
    .B1(_05404_),
    .B2(_05408_),
    .Y(_05409_)
  );
  sg13g2_nand2_1 _15387_ (
    .A(_03150_),
    .B(_07934_),
    .Y(_05410_)
  );
  sg13g2_o21ai_1 _15388_ (
    .A1(addr_i_3_),
    .A2(_03132_),
    .B1(_05410_),
    .Y(_05411_)
  );
  sg13g2_nand2_1 _15389_ (
    .A(_02437_),
    .B(_02742_),
    .Y(_05412_)
  );
  sg13g2_o21ai_1 _15390_ (
    .A1(_01231_),
    .A2(_02641_),
    .B1(_02344_),
    .Y(_05414_)
  );
  sg13g2_a21oi_1 _15391_ (
    .A1(_05412_),
    .A2(_05414_),
    .B1(_01911_),
    .Y(_05415_)
  );
  sg13g2_o21ai_1 _15392_ (
    .A1(_02107_),
    .A2(_08045_),
    .B1(addr_i_5_),
    .Y(_05416_)
  );
  sg13g2_o21ai_1 _15393_ (
    .A1(_00150_),
    .A2(_02501_),
    .B1(_05416_),
    .Y(_05417_)
  );
  sg13g2_a21oi_1 _15394_ (
    .A1(_05501_),
    .A2(_08045_),
    .B1(_01459_),
    .Y(_05418_)
  );
  sg13g2_o21ai_1 _15395_ (
    .A1(_00715_),
    .A2(_07879_),
    .B1(_08045_),
    .Y(_05419_)
  );
  sg13g2_o21ai_1 _15396_ (
    .A1(addr_i_3_),
    .A2(_05418_),
    .B1(_05419_),
    .Y(_05420_)
  );
  sg13g2_a21oi_1 _15397_ (
    .A1(addr_i_4_),
    .A2(_05417_),
    .B1(_05420_),
    .Y(_05421_)
  );
  sg13g2_a22oi_1 _15398_ (
    .A1(_00827_),
    .A2(_05411_),
    .B1(_05415_),
    .B2(_05421_),
    .Y(_05422_)
  );
  sg13g2_o21ai_1 _15399_ (
    .A1(addr_i_8_),
    .A2(_05409_),
    .B1(_05422_),
    .Y(_05423_)
  );
  sg13g2_nand2_1 _15400_ (
    .A(_00391_),
    .B(_01305_),
    .Y(_05425_)
  );
  sg13g2_a22oi_1 _15401_ (
    .A1(addr_i_3_),
    .A2(_05425_),
    .B1(_01845_),
    .B2(_00230_),
    .Y(_05426_)
  );
  sg13g2_nand2_1 _15402_ (
    .A(_07636_),
    .B(_09493_),
    .Y(_05427_)
  );
  sg13g2_o21ai_1 _15403_ (
    .A1(addr_i_4_),
    .A2(_03485_),
    .B1(_05427_),
    .Y(_05428_)
  );
  sg13g2_a21oi_1 _15404_ (
    .A1(_01077_),
    .A2(_03570_),
    .B1(addr_i_5_),
    .Y(_05429_)
  );
  sg13g2_nand2_1 _15405_ (
    .A(addr_i_2_),
    .B(_03875_),
    .Y(_05430_)
  );
  sg13g2_a21oi_1 _15406_ (
    .A1(_00140_),
    .A2(_05430_),
    .B1(_00554_),
    .Y(_05431_)
  );
  sg13g2_a22oi_1 _15407_ (
    .A1(_05867_),
    .A2(_05428_),
    .B1(_05429_),
    .B2(_05431_),
    .Y(_05432_)
  );
  sg13g2_nor2_1 _15408_ (
    .A(_06905_),
    .B(_05432_),
    .Y(_05433_)
  );
  sg13g2_a22oi_1 _15409_ (
    .A1(addr_i_3_),
    .A2(_03323_),
    .B1(_04098_),
    .B2(_00491_),
    .Y(_05434_)
  );
  sg13g2_o21ai_1 _15410_ (
    .A1(_00324_),
    .A2(_05434_),
    .B1(addr_i_8_),
    .Y(_05436_)
  );
  sg13g2_nor3_1 _15411_ (
    .A(_05426_),
    .B(_05433_),
    .C(_05436_),
    .Y(_05437_)
  );
  sg13g2_a21oi_1 _15412_ (
    .A1(_03424_),
    .A2(_07072_),
    .B1(_03854_),
    .Y(_05438_)
  );
  sg13g2_a21oi_1 _15413_ (
    .A1(addr_i_4_),
    .A2(_00582_),
    .B1(_03358_),
    .Y(_05439_)
  );
  sg13g2_nand2_1 _15414_ (
    .A(_05402_),
    .B(_02021_),
    .Y(_05440_)
  );
  sg13g2_a21oi_1 _15415_ (
    .A1(_01872_),
    .A2(_05440_),
    .B1(addr_i_7_),
    .Y(_05441_)
  );
  sg13g2_nor4_1 _15416_ (
    .A(addr_i_6_),
    .B(_05438_),
    .C(_05439_),
    .D(_05441_),
    .Y(_05442_)
  );
  sg13g2_nand3_1 _15417_ (
    .A(_00428_),
    .B(_00688_),
    .C(_01398_),
    .Y(_05443_)
  );
  sg13g2_a21oi_1 _15418_ (
    .A1(_00014_),
    .A2(_03665_),
    .B1(_08144_),
    .Y(_05444_)
  );
  sg13g2_o21ai_1 _15419_ (
    .A1(addr_i_3_),
    .A2(_01539_),
    .B1(_05444_),
    .Y(_05445_)
  );
  sg13g2_a21oi_1 _15420_ (
    .A1(_09486_),
    .A2(_05445_),
    .B1(addr_i_8_),
    .Y(_05447_)
  );
  sg13g2_o21ai_1 _15421_ (
    .A1(_01184_),
    .A2(_05443_),
    .B1(_05447_),
    .Y(_05448_)
  );
  sg13g2_o21ai_1 _15422_ (
    .A1(_05442_),
    .A2(_05448_),
    .B1(_01174_),
    .Y(_05449_)
  );
  sg13g2_o21ai_1 _15423_ (
    .A1(_05437_),
    .A2(_05449_),
    .B1(addr_i_11_),
    .Y(_05450_)
  );
  sg13g2_nand2_1 _15424_ (
    .A(_03953_),
    .B(_00620_),
    .Y(_05451_)
  );
  sg13g2_o21ai_1 _15425_ (
    .A1(_00199_),
    .A2(_01033_),
    .B1(addr_i_7_),
    .Y(_05452_)
  );
  sg13g2_a21oi_1 _15426_ (
    .A1(_00938_),
    .A2(_05452_),
    .B1(addr_i_2_),
    .Y(_05453_)
  );
  sg13g2_nand3_1 _15427_ (
    .A(_01113_),
    .B(_02053_),
    .C(_01384_),
    .Y(_05454_)
  );
  sg13g2_a21oi_1 _15428_ (
    .A1(_04087_),
    .A2(_05454_),
    .B1(addr_i_6_),
    .Y(_05455_)
  );
  sg13g2_a22oi_1 _15429_ (
    .A1(addr_i_4_),
    .A2(_05451_),
    .B1(_05453_),
    .B2(_05455_),
    .Y(_05456_)
  );
  sg13g2_o21ai_1 _15430_ (
    .A1(_06729_),
    .A2(_00242_),
    .B1(_01113_),
    .Y(_05458_)
  );
  sg13g2_nand3_1 _15431_ (
    .A(_04285_),
    .B(_08232_),
    .C(_05458_),
    .Y(_05459_)
  );
  sg13g2_nand2_1 _15432_ (
    .A(_01588_),
    .B(_00635_),
    .Y(_05460_)
  );
  sg13g2_a21oi_1 _15433_ (
    .A1(_00926_),
    .A2(_05460_),
    .B1(_00445_),
    .Y(_05461_)
  );
  sg13g2_a21oi_1 _15434_ (
    .A1(_00190_),
    .A2(_05459_),
    .B1(_05461_),
    .Y(_05462_)
  );
  sg13g2_o21ai_1 _15435_ (
    .A1(_00047_),
    .A2(_05456_),
    .B1(_05462_),
    .Y(_05463_)
  );
  sg13g2_nand2_1 _15436_ (
    .A(_02387_),
    .B(_02890_),
    .Y(_05464_)
  );
  sg13g2_nand4_1 _15437_ (
    .A(addr_i_7_),
    .B(_01224_),
    .C(_03131_),
    .D(_05464_),
    .Y(_05465_)
  );
  sg13g2_nor3_1 _15438_ (
    .A(_00479_),
    .B(_08288_),
    .C(_04225_),
    .Y(_05466_)
  );
  sg13g2_and2_1 _15439_ (
    .A(_02380_),
    .B(_04164_),
    .X(_05467_)
  );
  sg13g2_o21ai_1 _15440_ (
    .A1(_05466_),
    .A2(_05467_),
    .B1(_05218_),
    .Y(_05469_)
  );
  sg13g2_nor2_1 _15441_ (
    .A(_03267_),
    .B(_00177_),
    .Y(_05470_)
  );
  sg13g2_nand3_1 _15442_ (
    .A(addr_i_3_),
    .B(addr_i_7_),
    .C(_06862_),
    .Y(_05471_)
  );
  sg13g2_a21oi_1 _15443_ (
    .A1(_05470_),
    .A2(_05471_),
    .B1(addr_i_6_),
    .Y(_05472_)
  );
  sg13g2_a22oi_1 _15444_ (
    .A1(_05465_),
    .A2(_05469_),
    .B1(addr_i_8_),
    .B2(_05472_),
    .Y(_05473_)
  );
  sg13g2_a22oi_1 _15445_ (
    .A1(addr_i_8_),
    .A2(_05463_),
    .B1(_05473_),
    .B2(_01351_),
    .Y(_05474_)
  );
  sg13g2_a21oi_1 _15446_ (
    .A1(_00549_),
    .A2(_00566_),
    .B1(addr_i_3_),
    .Y(_05475_)
  );
  sg13g2_o21ai_1 _15447_ (
    .A1(_00342_),
    .A2(_02152_),
    .B1(addr_i_3_),
    .Y(_05476_)
  );
  sg13g2_a21oi_1 _15448_ (
    .A1(_03167_),
    .A2(_05476_),
    .B1(_08000_),
    .Y(_05477_)
  );
  sg13g2_a22oi_1 _15449_ (
    .A1(_02287_),
    .A2(_00568_),
    .B1(_05475_),
    .B2(_05477_),
    .Y(_05478_)
  );
  sg13g2_o21ai_1 _15450_ (
    .A1(addr_i_2_),
    .A2(_00299_),
    .B1(_02546_),
    .Y(_05480_)
  );
  sg13g2_o21ai_1 _15451_ (
    .A1(_07658_),
    .A2(_06220_),
    .B1(addr_i_7_),
    .Y(_05481_)
  );
  sg13g2_a21oi_1 _15452_ (
    .A1(_02815_),
    .A2(_05481_),
    .B1(addr_i_3_),
    .Y(_05482_)
  );
  sg13g2_a21oi_1 _15453_ (
    .A1(_03652_),
    .A2(_05480_),
    .B1(_05482_),
    .Y(_05483_)
  );
  sg13g2_o21ai_1 _15454_ (
    .A1(addr_i_7_),
    .A2(_05478_),
    .B1(_05483_),
    .Y(_05484_)
  );
  sg13g2_nand3_1 _15455_ (
    .A(addr_i_2_),
    .B(addr_i_5_),
    .C(_00025_),
    .Y(_05485_)
  );
  sg13g2_a21oi_1 _15456_ (
    .A1(_03540_),
    .A2(_05485_),
    .B1(addr_i_4_),
    .Y(_05486_)
  );
  sg13g2_o21ai_1 _15457_ (
    .A1(addr_i_2_),
    .A2(_02312_),
    .B1(_04640_),
    .Y(_05487_)
  );
  sg13g2_o21ai_1 _15458_ (
    .A1(_05486_),
    .A2(_05487_),
    .B1(addr_i_3_),
    .Y(_05488_)
  );
  sg13g2_xnor2_1 _15459_ (
    .A(_03908_),
    .B(_08597_),
    .Y(_05489_)
  );
  sg13g2_o21ai_1 _15460_ (
    .A1(_06729_),
    .A2(_03676_),
    .B1(addr_i_4_),
    .Y(_05491_)
  );
  sg13g2_o21ai_1 _15461_ (
    .A1(addr_i_6_),
    .A2(_05489_),
    .B1(_05491_),
    .Y(_05492_)
  );
  sg13g2_a21oi_1 _15462_ (
    .A1(_00726_),
    .A2(_05492_),
    .B1(_01604_),
    .Y(_05493_)
  );
  sg13g2_and3_1 _15463_ (
    .A(_03617_),
    .B(_05488_),
    .C(_05493_),
    .X(_05494_)
  );
  sg13g2_a22oi_1 _15464_ (
    .A1(addr_i_8_),
    .A2(_05484_),
    .B1(_05494_),
    .B2(addr_i_9_),
    .Y(_05495_)
  );
  sg13g2_nor3_1 _15465_ (
    .A(addr_i_10_),
    .B(_05474_),
    .C(_05495_),
    .Y(_05496_)
  );
  sg13g2_a22oi_1 _15466_ (
    .A1(_05214_),
    .A2(_05423_),
    .B1(_05450_),
    .B2(_05496_),
    .Y(_05497_)
  );
  sg13g2_o21ai_1 _15467_ (
    .A1(_02598_),
    .A2(_05568_),
    .B1(addr_i_3_),
    .Y(_05498_)
  );
  sg13g2_o21ai_1 _15468_ (
    .A1(_00467_),
    .A2(_00591_),
    .B1(_05498_),
    .Y(_05499_)
  );
  sg13g2_o21ai_1 _15469_ (
    .A1(_08653_),
    .A2(_00278_),
    .B1(_01528_),
    .Y(_05500_)
  );
  sg13g2_a21oi_1 _15470_ (
    .A1(_01144_),
    .A2(_05500_),
    .B1(addr_i_6_),
    .Y(_05503_)
  );
  sg13g2_o21ai_1 _15471_ (
    .A1(_05499_),
    .A2(_05503_),
    .B1(_06630_),
    .Y(_05504_)
  );
  sg13g2_o21ai_1 _15472_ (
    .A1(addr_i_2_),
    .A2(_02230_),
    .B1(_03559_),
    .Y(_05505_)
  );
  sg13g2_o21ai_1 _15473_ (
    .A1(_00269_),
    .A2(_02598_),
    .B1(_05402_),
    .Y(_05506_)
  );
  sg13g2_a21oi_1 _15474_ (
    .A1(_00339_),
    .A2(_05506_),
    .B1(_00485_),
    .Y(_05507_)
  );
  sg13g2_a22oi_1 _15475_ (
    .A1(addr_i_4_),
    .A2(_05505_),
    .B1(_05507_),
    .B2(_03520_),
    .Y(_05508_)
  );
  sg13g2_nor2_1 _15476_ (
    .A(addr_i_8_),
    .B(_05508_),
    .Y(_05509_)
  );
  sg13g2_nand3_1 _15477_ (
    .A(_00391_),
    .B(_01872_),
    .C(_05263_),
    .Y(_05510_)
  );
  sg13g2_o21ai_1 _15478_ (
    .A1(_00534_),
    .A2(_00947_),
    .B1(addr_i_4_),
    .Y(_05511_)
  );
  sg13g2_nor2_1 _15479_ (
    .A(_02602_),
    .B(_01276_),
    .Y(_05512_)
  );
  sg13g2_o21ai_1 _15480_ (
    .A1(_03577_),
    .A2(_05512_),
    .B1(_01674_),
    .Y(_05514_)
  );
  sg13g2_nand4_1 _15481_ (
    .A(_01354_),
    .B(_00478_),
    .C(_05511_),
    .D(_05514_),
    .Y(_05515_)
  );
  sg13g2_nand3_1 _15482_ (
    .A(addr_i_3_),
    .B(_00716_),
    .C(_01912_),
    .Y(_05516_)
  );
  sg13g2_o21ai_1 _15483_ (
    .A1(_07757_),
    .A2(_02424_),
    .B1(_01067_),
    .Y(_05517_)
  );
  sg13g2_nand3_1 _15484_ (
    .A(_01878_),
    .B(_05516_),
    .C(_05517_),
    .Y(_05518_)
  );
  sg13g2_nand2_1 _15485_ (
    .A(addr_i_8_),
    .B(_05518_),
    .Y(_05519_)
  );
  sg13g2_a221oi_1 _15486_ (
    .A1(_00402_),
    .A2(_05510_),
    .B1(_05515_),
    .B2(addr_i_7_),
    .C1(_05519_),
    .Y(_05520_)
  );
  sg13g2_a22oi_1 _15487_ (
    .A1(_05504_),
    .A2(_05509_),
    .B1(_06652_),
    .B2(_05520_),
    .Y(_05521_)
  );
  sg13g2_nor2_1 _15488_ (
    .A(_00825_),
    .B(_00270_),
    .Y(_05522_)
  );
  sg13g2_o21ai_1 _15489_ (
    .A1(_00070_),
    .A2(_06795_),
    .B1(_04296_),
    .Y(_05523_)
  );
  sg13g2_a21oi_1 _15490_ (
    .A1(_00951_),
    .A2(_02573_),
    .B1(_01125_),
    .Y(_05525_)
  );
  sg13g2_a22oi_1 _15491_ (
    .A1(_07149_),
    .A2(_05523_),
    .B1(_05525_),
    .B2(addr_i_6_),
    .Y(_05526_)
  );
  sg13g2_o21ai_1 _15492_ (
    .A1(_00258_),
    .A2(_02241_),
    .B1(_05600_),
    .Y(_05527_)
  );
  sg13g2_nand2_1 _15493_ (
    .A(addr_i_8_),
    .B(_05527_),
    .Y(_05528_)
  );
  sg13g2_a22oi_1 _15494_ (
    .A1(_04156_),
    .A2(_05522_),
    .B1(_05526_),
    .B2(_05528_),
    .Y(_05529_)
  );
  sg13g2_nor3_1 _15495_ (
    .A(_02759_),
    .B(_00279_),
    .C(_05195_),
    .Y(_05530_)
  );
  sg13g2_nor4_1 _15496_ (
    .A(_00492_),
    .B(_05568_),
    .C(_01246_),
    .D(_04490_),
    .Y(_05531_)
  );
  sg13g2_nand3_1 _15497_ (
    .A(_05218_),
    .B(_00762_),
    .C(_05479_),
    .Y(_05532_)
  );
  sg13g2_o21ai_1 _15498_ (
    .A1(_08343_),
    .A2(_09083_),
    .B1(addr_i_3_),
    .Y(_05533_)
  );
  sg13g2_nand3_1 _15499_ (
    .A(addr_i_7_),
    .B(_00651_),
    .C(_05533_),
    .Y(_05534_)
  );
  sg13g2_a21oi_1 _15500_ (
    .A1(_05532_),
    .A2(_05534_),
    .B1(addr_i_6_),
    .Y(_05536_)
  );
  sg13g2_nor4_1 _15501_ (
    .A(addr_i_8_),
    .B(_05530_),
    .C(_05531_),
    .D(_05536_),
    .Y(_05537_)
  );
  sg13g2_nor3_1 _15502_ (
    .A(_00925_),
    .B(_05529_),
    .C(_05537_),
    .Y(_05538_)
  );
  sg13g2_nand2_1 _15503_ (
    .A(addr_i_3_),
    .B(_03905_),
    .Y(_05539_)
  );
  sg13g2_o21ai_1 _15504_ (
    .A1(_06176_),
    .A2(_04265_),
    .B1(addr_i_4_),
    .Y(_05540_)
  );
  sg13g2_a21oi_1 _15505_ (
    .A1(_05539_),
    .A2(_05540_),
    .B1(addr_i_7_),
    .Y(_05541_)
  );
  sg13g2_o21ai_1 _15506_ (
    .A1(addr_i_4_),
    .A2(_02108_),
    .B1(_04793_),
    .Y(_05542_)
  );
  sg13g2_nand2b_1 _15507_ (
    .A_N(_05542_),
    .B(addr_i_2_),
    .Y(_05543_)
  );
  sg13g2_nor2_1 _15508_ (
    .A(addr_i_3_),
    .B(_01461_),
    .Y(_05544_)
  );
  sg13g2_a221oi_1 _15509_ (
    .A1(_04060_),
    .A2(_05543_),
    .B1(_05544_),
    .B2(_00148_),
    .C1(_02064_),
    .Y(_05545_)
  );
  sg13g2_o21ai_1 _15510_ (
    .A1(_01867_),
    .A2(_06563_),
    .B1(_08166_),
    .Y(_05547_)
  );
  sg13g2_a21oi_1 _15511_ (
    .A1(_02695_),
    .A2(_05547_),
    .B1(addr_i_3_),
    .Y(_05548_)
  );
  sg13g2_o21ai_1 _15512_ (
    .A1(_00138_),
    .A2(_08951_),
    .B1(addr_i_8_),
    .Y(_05549_)
  );
  sg13g2_nor4_1 _15513_ (
    .A(_05541_),
    .B(_05545_),
    .C(_05548_),
    .D(_05549_),
    .Y(_05550_)
  );
  sg13g2_o21ai_1 _15514_ (
    .A1(addr_i_7_),
    .A2(_03172_),
    .B1(_00120_),
    .Y(_05551_)
  );
  sg13g2_a21oi_1 _15515_ (
    .A1(_01791_),
    .A2(_05551_),
    .B1(_01970_),
    .Y(_05552_)
  );
  sg13g2_o21ai_1 _15516_ (
    .A1(_00732_),
    .A2(_05552_),
    .B1(addr_i_4_),
    .Y(_05553_)
  );
  sg13g2_o21ai_1 _15517_ (
    .A1(addr_i_5_),
    .A2(_07812_),
    .B1(_07359_),
    .Y(_05554_)
  );
  sg13g2_nor2_1 _15518_ (
    .A(_08044_),
    .B(_00664_),
    .Y(_05555_)
  );
  sg13g2_a22oi_1 _15519_ (
    .A1(addr_i_3_),
    .A2(_05555_),
    .B1(_02119_),
    .B2(addr_i_7_),
    .Y(_05556_)
  );
  sg13g2_nand2_1 _15520_ (
    .A(_01077_),
    .B(_00571_),
    .Y(_05558_)
  );
  sg13g2_nor2_1 _15521_ (
    .A(_09149_),
    .B(_05558_),
    .Y(_05559_)
  );
  sg13g2_a22oi_1 _15522_ (
    .A1(_05554_),
    .A2(_05556_),
    .B1(_05559_),
    .B2(addr_i_8_),
    .Y(_05560_)
  );
  sg13g2_a21oi_1 _15523_ (
    .A1(_05553_),
    .A2(_05560_),
    .B1(addr_i_9_),
    .Y(_05561_)
  );
  sg13g2_nand2b_1 _15524_ (
    .A_N(_05550_),
    .B(_05561_),
    .Y(_05562_)
  );
  sg13g2_nor2_1 _15525_ (
    .A(_02645_),
    .B(_05036_),
    .Y(_05563_)
  );
  sg13g2_o21ai_1 _15526_ (
    .A1(_04957_),
    .A2(_05563_),
    .B1(_05070_),
    .Y(_05564_)
  );
  sg13g2_a21oi_1 _15527_ (
    .A1(_04362_),
    .A2(_00019_),
    .B1(_00961_),
    .Y(_05565_)
  );
  sg13g2_nor2_1 _15528_ (
    .A(_01910_),
    .B(_05565_),
    .Y(_05566_)
  );
  sg13g2_a21o_1 _15529_ (
    .A1(_05564_),
    .A2(_05566_),
    .B1(_00091_),
    .X(_05567_)
  );
  sg13g2_nand2_1 _15530_ (
    .A(addr_i_3_),
    .B(_05003_),
    .Y(_05569_)
  );
  sg13g2_nand3_1 _15531_ (
    .A(_00262_),
    .B(_00458_),
    .C(_05569_),
    .Y(_05570_)
  );
  sg13g2_nand3_1 _15532_ (
    .A(_09473_),
    .B(_00871_),
    .C(_05334_),
    .Y(_05571_)
  );
  sg13g2_nand4_1 _15533_ (
    .A(addr_i_8_),
    .B(_05567_),
    .C(_05570_),
    .D(_05571_),
    .Y(_05572_)
  );
  sg13g2_o21ai_1 _15534_ (
    .A1(addr_i_3_),
    .A2(_00154_),
    .B1(_00246_),
    .Y(_05573_)
  );
  sg13g2_o21ai_1 _15535_ (
    .A1(_00977_),
    .A2(_05573_),
    .B1(addr_i_4_),
    .Y(_05574_)
  );
  sg13g2_nor2_1 _15536_ (
    .A(addr_i_4_),
    .B(_03413_),
    .Y(_05575_)
  );
  sg13g2_o21ai_1 _15537_ (
    .A1(_05575_),
    .A2(_00226_),
    .B1(addr_i_3_),
    .Y(_05576_)
  );
  sg13g2_a21oi_1 _15538_ (
    .A1(_05574_),
    .A2(_05576_),
    .B1(addr_i_6_),
    .Y(_05577_)
  );
  sg13g2_o21ai_1 _15539_ (
    .A1(_00117_),
    .A2(_00608_),
    .B1(_01120_),
    .Y(_05578_)
  );
  sg13g2_o21ai_1 _15540_ (
    .A1(addr_i_3_),
    .A2(_03905_),
    .B1(_00019_),
    .Y(_05580_)
  );
  sg13g2_a22oi_1 _15541_ (
    .A1(_01120_),
    .A2(_05580_),
    .B1(_02598_),
    .B2(addr_i_7_),
    .Y(_05581_)
  );
  sg13g2_a21oi_1 _15542_ (
    .A1(_04246_),
    .A2(_05578_),
    .B1(_05581_),
    .Y(_05582_)
  );
  sg13g2_or3_1 _15543_ (
    .A(addr_i_8_),
    .B(_05577_),
    .C(_05582_),
    .X(_05583_)
  );
  sg13g2_nand3_1 _15544_ (
    .A(addr_i_9_),
    .B(_05572_),
    .C(_05583_),
    .Y(_05584_)
  );
  sg13g2_a21oi_1 _15545_ (
    .A1(_05562_),
    .A2(_05584_),
    .B1(addr_i_10_),
    .Y(_05585_)
  );
  sg13g2_nor4_1 _15546_ (
    .A(addr_i_11_),
    .B(_05521_),
    .C(_05538_),
    .D(_05585_),
    .Y(_05586_)
  );
  sg13g2_or3_1 _15547_ (
    .A(addr_i_12_),
    .B(_05497_),
    .C(_05586_),
    .X(_05587_)
  );
  sg13g2_o21ai_1 _15548_ (
    .A1(_02251_),
    .A2(_05399_),
    .B1(_05587_),
    .Y(data_o_24_)
  );
  sg13g2_nor2_1 _15549_ (
    .A(_02569_),
    .B(_00719_),
    .Y(_05588_)
  );
  sg13g2_nor2_1 _15550_ (
    .A(_03798_),
    .B(_03875_),
    .Y(_05590_)
  );
  sg13g2_a21oi_1 _15551_ (
    .A1(addr_i_3_),
    .A2(_02080_),
    .B1(_05590_),
    .Y(_05591_)
  );
  sg13g2_nor2_1 _15552_ (
    .A(addr_i_2_),
    .B(_05591_),
    .Y(_05592_)
  );
  sg13g2_o21ai_1 _15553_ (
    .A1(_05588_),
    .A2(_05592_),
    .B1(_01630_),
    .Y(_05593_)
  );
  sg13g2_a22oi_1 _15554_ (
    .A1(_09127_),
    .A2(_07248_),
    .B1(_00644_),
    .B2(_08752_),
    .Y(_05594_)
  );
  sg13g2_nor3_1 _15555_ (
    .A(addr_i_3_),
    .B(_02265_),
    .C(_05932_),
    .Y(_05595_)
  );
  sg13g2_nand2_1 _15556_ (
    .A(addr_i_4_),
    .B(_00454_),
    .Y(_05596_)
  );
  sg13g2_o21ai_1 _15557_ (
    .A1(_05594_),
    .A2(_05595_),
    .B1(_05596_),
    .Y(_05597_)
  );
  sg13g2_o21ai_1 _15558_ (
    .A1(_03431_),
    .A2(_00825_),
    .B1(addr_i_8_),
    .Y(_05598_)
  );
  sg13g2_nand2_1 _15559_ (
    .A(addr_i_3_),
    .B(_05280_),
    .Y(_05599_)
  );
  sg13g2_a21oi_1 _15560_ (
    .A1(_00069_),
    .A2(_05599_),
    .B1(_02513_),
    .Y(_05601_)
  );
  sg13g2_a22oi_1 _15561_ (
    .A1(addr_i_2_),
    .A2(_05597_),
    .B1(_05598_),
    .B2(_05601_),
    .Y(_05602_)
  );
  sg13g2_nor2_1 _15562_ (
    .A(addr_i_4_),
    .B(_08376_),
    .Y(_05603_)
  );
  sg13g2_a21oi_1 _15563_ (
    .A1(addr_i_5_),
    .A2(_08929_),
    .B1(_00484_),
    .Y(_05604_)
  );
  sg13g2_o21ai_1 _15564_ (
    .A1(_05603_),
    .A2(_05604_),
    .B1(_04461_),
    .Y(_05605_)
  );
  sg13g2_o21ai_1 _15565_ (
    .A1(_00070_),
    .A2(_02954_),
    .B1(_05605_),
    .Y(_05606_)
  );
  sg13g2_o21ai_1 _15566_ (
    .A1(addr_i_5_),
    .A2(_03690_),
    .B1(addr_i_3_),
    .Y(_05607_)
  );
  sg13g2_a21oi_1 _15567_ (
    .A1(_00484_),
    .A2(_08254_),
    .B1(_09509_),
    .Y(_05608_)
  );
  sg13g2_a21oi_1 _15568_ (
    .A1(_00554_),
    .A2(_01718_),
    .B1(_05608_),
    .Y(_05609_)
  );
  sg13g2_a21oi_1 _15569_ (
    .A1(_05607_),
    .A2(_05609_),
    .B1(addr_i_2_),
    .Y(_05610_)
  );
  sg13g2_nand2_1 _15570_ (
    .A(_00104_),
    .B(_08520_),
    .Y(_05613_)
  );
  sg13g2_a21oi_1 _15571_ (
    .A1(addr_i_3_),
    .A2(_05613_),
    .B1(_02265_),
    .Y(_05614_)
  );
  sg13g2_o21ai_1 _15572_ (
    .A1(addr_i_7_),
    .A2(_05614_),
    .B1(_00943_),
    .Y(_05615_)
  );
  sg13g2_a22oi_1 _15573_ (
    .A1(addr_i_2_),
    .A2(_05606_),
    .B1(_05610_),
    .B2(_05615_),
    .Y(_05616_)
  );
  sg13g2_nor2_1 _15574_ (
    .A(addr_i_8_),
    .B(_05616_),
    .Y(_05617_)
  );
  sg13g2_a22oi_1 _15575_ (
    .A1(_05593_),
    .A2(_05602_),
    .B1(_05617_),
    .B2(_09326_),
    .Y(_05618_)
  );
  sg13g2_o21ai_1 _15576_ (
    .A1(addr_i_4_),
    .A2(_05833_),
    .B1(_06784_),
    .Y(_05619_)
  );
  sg13g2_a21oi_1 _15577_ (
    .A1(_02191_),
    .A2(_01441_),
    .B1(_04251_),
    .Y(_05620_)
  );
  sg13g2_o21ai_1 _15578_ (
    .A1(_02513_),
    .A2(_00760_),
    .B1(_04296_),
    .Y(_05621_)
  );
  sg13g2_a22oi_1 _15579_ (
    .A1(addr_i_2_),
    .A2(_05619_),
    .B1(_05620_),
    .B2(_05621_),
    .Y(_05622_)
  );
  sg13g2_a21oi_1 _15580_ (
    .A1(addr_i_2_),
    .A2(_00275_),
    .B1(_00158_),
    .Y(_05624_)
  );
  sg13g2_o21ai_1 _15581_ (
    .A1(_01114_),
    .A2(_05624_),
    .B1(_01212_),
    .Y(_05625_)
  );
  sg13g2_a21oi_1 _15582_ (
    .A1(_01543_),
    .A2(_04916_),
    .B1(addr_i_4_),
    .Y(_05626_)
  );
  sg13g2_a22oi_1 _15583_ (
    .A1(_01935_),
    .A2(_05625_),
    .B1(_05626_),
    .B2(_04499_),
    .Y(_05627_)
  );
  sg13g2_o21ai_1 _15584_ (
    .A1(_00191_),
    .A2(_05622_),
    .B1(_05627_),
    .Y(_05628_)
  );
  sg13g2_a21oi_1 _15585_ (
    .A1(_02371_),
    .A2(_02283_),
    .B1(addr_i_4_),
    .Y(_05629_)
  );
  sg13g2_a21o_1 _15586_ (
    .A1(addr_i_4_),
    .A2(_04572_),
    .B1(_05629_),
    .X(_05630_)
  );
  sg13g2_nor2_1 _15587_ (
    .A(_02294_),
    .B(_01001_),
    .Y(_05631_)
  );
  sg13g2_a221oi_1 _15588_ (
    .A1(_01215_),
    .A2(_04048_),
    .B1(_05630_),
    .B2(addr_i_2_),
    .C1(_05631_),
    .Y(_05632_)
  );
  sg13g2_a21oi_1 _15589_ (
    .A1(_00482_),
    .A2(_02048_),
    .B1(addr_i_7_),
    .Y(_05633_)
  );
  sg13g2_nor3_1 _15590_ (
    .A(addr_i_3_),
    .B(_02772_),
    .C(_05633_),
    .Y(_05635_)
  );
  sg13g2_a21oi_1 _15591_ (
    .A1(addr_i_3_),
    .A2(_05632_),
    .B1(_05635_),
    .Y(_05636_)
  );
  sg13g2_nor3_1 _15592_ (
    .A(addr_i_8_),
    .B(_04506_),
    .C(_05636_),
    .Y(_05637_)
  );
  sg13g2_a22oi_1 _15593_ (
    .A1(addr_i_8_),
    .A2(_05628_),
    .B1(_05637_),
    .B2(addr_i_9_),
    .Y(_05638_)
  );
  sg13g2_nor2_1 _15594_ (
    .A(addr_i_11_),
    .B(_03841_),
    .Y(_05639_)
  );
  sg13g2_o21ai_1 _15595_ (
    .A1(_05618_),
    .A2(_05638_),
    .B1(_05639_),
    .Y(_05640_)
  );
  sg13g2_o21ai_1 _15596_ (
    .A1(addr_i_3_),
    .A2(_00901_),
    .B1(_07337_),
    .Y(_05641_)
  );
  sg13g2_o21ai_1 _15597_ (
    .A1(_00531_),
    .A2(_03089_),
    .B1(_01518_),
    .Y(_05642_)
  );
  sg13g2_a21oi_1 _15598_ (
    .A1(_09476_),
    .A2(_00820_),
    .B1(addr_i_6_),
    .Y(_05643_)
  );
  sg13g2_a22oi_1 _15599_ (
    .A1(addr_i_4_),
    .A2(_05641_),
    .B1(_05642_),
    .B2(_05643_),
    .Y(_05644_)
  );
  sg13g2_nor3_1 _15600_ (
    .A(_00261_),
    .B(_00999_),
    .C(_08807_),
    .Y(_05646_)
  );
  sg13g2_o21ai_1 _15601_ (
    .A1(_03793_),
    .A2(_05646_),
    .B1(addr_i_4_),
    .Y(_05647_)
  );
  sg13g2_nand2_1 _15602_ (
    .A(_04749_),
    .B(_01943_),
    .Y(_05648_)
  );
  sg13g2_a21oi_1 _15603_ (
    .A1(_08266_),
    .A2(_05648_),
    .B1(addr_i_4_),
    .Y(_05649_)
  );
  sg13g2_a22oi_1 _15604_ (
    .A1(addr_i_3_),
    .A2(_00128_),
    .B1(_00600_),
    .B2(_05649_),
    .Y(_05650_)
  );
  sg13g2_a21oi_1 _15605_ (
    .A1(addr_i_4_),
    .A2(addr_i_5_),
    .B1(addr_i_6_),
    .Y(_05651_)
  );
  sg13g2_inv_1 _15606_ (
    .A(_05651_),
    .Y(_05652_)
  );
  sg13g2_a21oi_1 _15607_ (
    .A1(_01067_),
    .A2(_05652_),
    .B1(_01436_),
    .Y(_05653_)
  );
  sg13g2_o21ai_1 _15608_ (
    .A1(addr_i_2_),
    .A2(_05653_),
    .B1(_00185_),
    .Y(_05654_)
  );
  sg13g2_a21oi_1 _15609_ (
    .A1(_00567_),
    .A2(_02822_),
    .B1(_00315_),
    .Y(_05655_)
  );
  sg13g2_a22oi_1 _15610_ (
    .A1(_06905_),
    .A2(_05654_),
    .B1(_05655_),
    .B2(_03975_),
    .Y(_05657_)
  );
  sg13g2_a21oi_1 _15611_ (
    .A1(_05647_),
    .A2(_05650_),
    .B1(_05657_),
    .Y(_05658_)
  );
  sg13g2_nor3_1 _15612_ (
    .A(_02700_),
    .B(_04152_),
    .C(_03030_),
    .Y(_05659_)
  );
  sg13g2_a21oi_1 _15613_ (
    .A1(_09326_),
    .A2(_05658_),
    .B1(_05659_),
    .Y(_05660_)
  );
  sg13g2_nor2_1 _15614_ (
    .A(_03040_),
    .B(addr_i_10_),
    .Y(_05661_)
  );
  sg13g2_o21ai_1 _15615_ (
    .A1(_05644_),
    .A2(_05660_),
    .B1(_05661_),
    .Y(_05662_)
  );
  sg13g2_o21ai_1 _15616_ (
    .A1(_01041_),
    .A2(_03287_),
    .B1(addr_i_6_),
    .Y(_05663_)
  );
  sg13g2_nand2_1 _15617_ (
    .A(_06784_),
    .B(_03457_),
    .Y(_05664_)
  );
  sg13g2_a22oi_1 _15618_ (
    .A1(addr_i_4_),
    .A2(_05664_),
    .B1(_05590_),
    .B2(_02203_),
    .Y(_05665_)
  );
  sg13g2_nand2b_1 _15619_ (
    .A_N(_05665_),
    .B(addr_i_2_),
    .Y(_05666_)
  );
  sg13g2_nand3_1 _15620_ (
    .A(_00047_),
    .B(addr_i_7_),
    .C(_00118_),
    .Y(_05668_)
  );
  sg13g2_nand3_1 _15621_ (
    .A(addr_i_3_),
    .B(_00292_),
    .C(_05542_),
    .Y(_05669_)
  );
  sg13g2_nand4_1 _15622_ (
    .A(_05663_),
    .B(_05666_),
    .C(_05668_),
    .D(_05669_),
    .Y(_05670_)
  );
  sg13g2_nand2_1 _15623_ (
    .A(_07503_),
    .B(_02103_),
    .Y(_05671_)
  );
  sg13g2_o21ai_1 _15624_ (
    .A1(_00103_),
    .A2(_00688_),
    .B1(_05671_),
    .Y(_05672_)
  );
  sg13g2_a21oi_1 _15625_ (
    .A1(_00072_),
    .A2(_01672_),
    .B1(_01194_),
    .Y(_05673_)
  );
  sg13g2_o21ai_1 _15626_ (
    .A1(_05280_),
    .A2(_07879_),
    .B1(addr_i_2_),
    .Y(_05674_)
  );
  sg13g2_nand3_1 _15627_ (
    .A(addr_i_6_),
    .B(_05673_),
    .C(_05674_),
    .Y(_05675_)
  );
  sg13g2_o21ai_1 _15628_ (
    .A1(addr_i_6_),
    .A2(_05672_),
    .B1(_05675_),
    .Y(_05676_)
  );
  sg13g2_o21ai_1 _15629_ (
    .A1(_02154_),
    .A2(_01567_),
    .B1(addr_i_3_),
    .Y(_05677_)
  );
  sg13g2_a21oi_1 _15630_ (
    .A1(_05676_),
    .A2(_05677_),
    .B1(addr_i_8_),
    .Y(_05679_)
  );
  sg13g2_a22oi_1 _15631_ (
    .A1(addr_i_8_),
    .A2(_05670_),
    .B1(_05679_),
    .B2(_09326_),
    .Y(_05680_)
  );
  sg13g2_a22oi_1 _15632_ (
    .A1(addr_i_2_),
    .A2(_04426_),
    .B1(_00569_),
    .B2(_00825_),
    .Y(_05681_)
  );
  sg13g2_a21oi_1 _15633_ (
    .A1(_02578_),
    .A2(_00712_),
    .B1(_00899_),
    .Y(_05682_)
  );
  sg13g2_nor3_1 _15634_ (
    .A(_05711_),
    .B(_03245_),
    .C(_07359_),
    .Y(_05683_)
  );
  sg13g2_o21ai_1 _15635_ (
    .A1(_06574_),
    .A2(_05683_),
    .B1(addr_i_5_),
    .Y(_05684_)
  );
  sg13g2_o21ai_1 _15636_ (
    .A1(_01024_),
    .A2(_03455_),
    .B1(_00799_),
    .Y(_05685_)
  );
  sg13g2_a21oi_1 _15637_ (
    .A1(_05684_),
    .A2(_05685_),
    .B1(addr_i_7_),
    .Y(_05686_)
  );
  sg13g2_nor4_1 _15638_ (
    .A(_00214_),
    .B(_05681_),
    .C(_05682_),
    .D(_05686_),
    .Y(_05687_)
  );
  sg13g2_a21oi_1 _15639_ (
    .A1(_02744_),
    .A2(_00430_),
    .B1(_00666_),
    .Y(_05688_)
  );
  sg13g2_a22oi_1 _15640_ (
    .A1(_01169_),
    .A2(_01716_),
    .B1(_02774_),
    .B2(_05688_),
    .Y(_05690_)
  );
  sg13g2_nor2_1 _15641_ (
    .A(_00779_),
    .B(_05690_),
    .Y(_05691_)
  );
  sg13g2_o21ai_1 _15642_ (
    .A1(_02105_),
    .A2(_03089_),
    .B1(_02807_),
    .Y(_05692_)
  );
  sg13g2_a22oi_1 _15643_ (
    .A1(addr_i_3_),
    .A2(_02943_),
    .B1(_03833_),
    .B2(_01155_),
    .Y(_05693_)
  );
  sg13g2_a22oi_1 _15644_ (
    .A1(_05600_),
    .A2(_05692_),
    .B1(_05693_),
    .B2(_01611_),
    .Y(_05694_)
  );
  sg13g2_nor2b_1 _15645_ (
    .A(_05691_),
    .B_N(_05694_),
    .Y(_05695_)
  );
  sg13g2_nor4_1 _15646_ (
    .A(addr_i_11_),
    .B(addr_i_10_),
    .C(_05687_),
    .D(_05695_),
    .Y(_05696_)
  );
  sg13g2_nand2b_1 _15647_ (
    .A_N(_05680_),
    .B(_05696_),
    .Y(_05697_)
  );
  sg13g2_o21ai_1 _15648_ (
    .A1(_06398_),
    .A2(_05932_),
    .B1(_06054_),
    .Y(_05698_)
  );
  sg13g2_a21oi_1 _15649_ (
    .A1(_07547_),
    .A2(_00542_),
    .B1(_06630_),
    .Y(_05699_)
  );
  sg13g2_nand2_1 _15650_ (
    .A(_05698_),
    .B(_05699_),
    .Y(_05701_)
  );
  sg13g2_nand4_1 _15651_ (
    .A(addr_i_4_),
    .B(addr_i_11_),
    .C(_01350_),
    .D(_05701_),
    .Y(_05702_)
  );
  sg13g2_nand4_1 _15652_ (
    .A(_05640_),
    .B(_05662_),
    .C(_05697_),
    .D(_05702_),
    .Y(_05703_)
  );
  sg13g2_o21ai_1 _15653_ (
    .A1(_00465_),
    .A2(_01376_),
    .B1(_01382_),
    .Y(_05704_)
  );
  sg13g2_a21oi_1 _15654_ (
    .A1(_08431_),
    .A2(_01060_),
    .B1(_01520_),
    .Y(_05705_)
  );
  sg13g2_o21ai_1 _15655_ (
    .A1(addr_i_3_),
    .A2(_07248_),
    .B1(_02287_),
    .Y(_05706_)
  );
  sg13g2_a21oi_1 _15656_ (
    .A1(_01104_),
    .A2(_05706_),
    .B1(addr_i_6_),
    .Y(_05707_)
  );
  sg13g2_o21ai_1 _15657_ (
    .A1(_05705_),
    .A2(_05707_),
    .B1(_00610_),
    .Y(_05708_)
  );
  sg13g2_a21oi_1 _15658_ (
    .A1(_00155_),
    .A2(_02683_),
    .B1(_04461_),
    .Y(_05709_)
  );
  sg13g2_nand2_1 _15659_ (
    .A(_04450_),
    .B(_05036_),
    .Y(_05710_)
  );
  sg13g2_a21oi_1 _15660_ (
    .A1(_01473_),
    .A2(_05710_),
    .B1(addr_i_6_),
    .Y(_05712_)
  );
  sg13g2_nor4_1 _15661_ (
    .A(_05568_),
    .B(_01285_),
    .C(_05709_),
    .D(_05712_),
    .Y(_05713_)
  );
  sg13g2_a22oi_1 _15662_ (
    .A1(addr_i_5_),
    .A2(_01339_),
    .B1(_00151_),
    .B2(_00600_),
    .Y(_05714_)
  );
  sg13g2_a21oi_1 _15663_ (
    .A1(_00831_),
    .A2(_00884_),
    .B1(_03132_),
    .Y(_05715_)
  );
  sg13g2_o21ai_1 _15664_ (
    .A1(_01380_),
    .A2(_00494_),
    .B1(_02501_),
    .Y(_05716_)
  );
  sg13g2_nand2b_1 _15665_ (
    .A_N(_05715_),
    .B(_05716_),
    .Y(_05717_)
  );
  sg13g2_nor3_1 _15666_ (
    .A(_05713_),
    .B(_05714_),
    .C(_05717_),
    .Y(_05718_)
  );
  sg13g2_nand3_1 _15667_ (
    .A(_05704_),
    .B(_05708_),
    .C(_05718_),
    .Y(_05719_)
  );
  sg13g2_nand2b_1 _15668_ (
    .A_N(_01305_),
    .B(_00822_),
    .Y(_05720_)
  );
  sg13g2_a21oi_1 _15669_ (
    .A1(_01108_),
    .A2(_05720_),
    .B1(addr_i_7_),
    .Y(_05721_)
  );
  sg13g2_a21oi_1 _15670_ (
    .A1(addr_i_3_),
    .A2(_03129_),
    .B1(_03033_),
    .Y(_05724_)
  );
  sg13g2_o21ai_1 _15671_ (
    .A1(_05822_),
    .A2(_05724_),
    .B1(_06508_),
    .Y(_05725_)
  );
  sg13g2_o21ai_1 _15672_ (
    .A1(_05721_),
    .A2(_05725_),
    .B1(addr_i_6_),
    .Y(_05726_)
  );
  sg13g2_o21ai_1 _15673_ (
    .A1(_00503_),
    .A2(_03012_),
    .B1(addr_i_4_),
    .Y(_05727_)
  );
  sg13g2_a21oi_1 _15674_ (
    .A1(_00999_),
    .A2(_04355_),
    .B1(_03455_),
    .Y(_05728_)
  );
  sg13g2_nand2_1 _15675_ (
    .A(_05727_),
    .B(_05728_),
    .Y(_05729_)
  );
  sg13g2_a21oi_1 _15676_ (
    .A1(addr_i_7_),
    .A2(_05729_),
    .B1(_02391_),
    .Y(_05730_)
  );
  sg13g2_a21oi_1 _15677_ (
    .A1(_05726_),
    .A2(_05730_),
    .B1(_02368_),
    .Y(_05731_)
  );
  sg13g2_o21ai_1 _15678_ (
    .A1(addr_i_7_),
    .A2(_02462_),
    .B1(addr_i_4_),
    .Y(_05732_)
  );
  sg13g2_a21oi_1 _15679_ (
    .A1(_00695_),
    .A2(_05732_),
    .B1(addr_i_2_),
    .Y(_05733_)
  );
  sg13g2_a21oi_1 _15680_ (
    .A1(_01615_),
    .A2(_02930_),
    .B1(addr_i_3_),
    .Y(_05735_)
  );
  sg13g2_o21ai_1 _15681_ (
    .A1(_05733_),
    .A2(_05735_),
    .B1(_01324_),
    .Y(_05736_)
  );
  sg13g2_nor2_1 _15682_ (
    .A(addr_i_7_),
    .B(_00304_),
    .Y(_05737_)
  );
  sg13g2_a21oi_1 _15683_ (
    .A1(_03820_),
    .A2(_01160_),
    .B1(addr_i_3_),
    .Y(_05738_)
  );
  sg13g2_nand2_1 _15684_ (
    .A(addr_i_5_),
    .B(_02529_),
    .Y(_05739_)
  );
  sg13g2_a22oi_1 _15685_ (
    .A1(_00305_),
    .A2(_00789_),
    .B1(_05738_),
    .B2(_05739_),
    .Y(_05740_)
  );
  sg13g2_a22oi_1 _15686_ (
    .A1(_00542_),
    .A2(_05737_),
    .B1(_05740_),
    .B2(_01611_),
    .Y(_05741_)
  );
  sg13g2_a21o_1 _15687_ (
    .A1(_05736_),
    .A2(_05741_),
    .B1(_01773_),
    .X(_05742_)
  );
  sg13g2_a22oi_1 _15688_ (
    .A1(addr_i_9_),
    .A2(_05719_),
    .B1(_05731_),
    .B2(_05742_),
    .Y(_05743_)
  );
  sg13g2_nor3_1 _15689_ (
    .A(_00015_),
    .B(_07945_),
    .C(_01846_),
    .Y(_05744_)
  );
  sg13g2_xor2_1 _15690_ (
    .A(addr_i_3_),
    .B(addr_i_5_),
    .X(_05746_)
  );
  sg13g2_xnor2_1 _15691_ (
    .A(_00408_),
    .B(_05746_),
    .Y(_05747_)
  );
  sg13g2_o21ai_1 _15692_ (
    .A1(_08045_),
    .A2(_05747_),
    .B1(_00385_),
    .Y(_05748_)
  );
  sg13g2_nand2_1 _15693_ (
    .A(_00339_),
    .B(_00704_),
    .Y(_05749_)
  );
  sg13g2_nor2_1 _15694_ (
    .A(_07425_),
    .B(_07668_),
    .Y(_05750_)
  );
  sg13g2_a22oi_1 _15695_ (
    .A1(_05258_),
    .A2(_03864_),
    .B1(_06497_),
    .B2(addr_i_4_),
    .Y(_05751_)
  );
  sg13g2_a21oi_1 _15696_ (
    .A1(addr_i_4_),
    .A2(_05750_),
    .B1(_05751_),
    .Y(_05752_)
  );
  sg13g2_a22oi_1 _15697_ (
    .A1(_04052_),
    .A2(_05749_),
    .B1(_05752_),
    .B2(_07614_),
    .Y(_05753_)
  );
  sg13g2_a22oi_1 _15698_ (
    .A1(_00884_),
    .A2(_05744_),
    .B1(_05748_),
    .B2(_05753_),
    .Y(_05754_)
  );
  sg13g2_a22oi_1 _15699_ (
    .A1(addr_i_4_),
    .A2(_01179_),
    .B1(_03501_),
    .B2(_06276_),
    .Y(_05755_)
  );
  sg13g2_nand2_1 _15700_ (
    .A(_01581_),
    .B(_00591_),
    .Y(_05757_)
  );
  sg13g2_a21oi_1 _15701_ (
    .A1(_00967_),
    .A2(_05757_),
    .B1(addr_i_3_),
    .Y(_05758_)
  );
  sg13g2_a22oi_1 _15702_ (
    .A1(addr_i_3_),
    .A2(_05755_),
    .B1(_05758_),
    .B2(_08830_),
    .Y(_05759_)
  );
  sg13g2_o21ai_1 _15703_ (
    .A1(_00824_),
    .A2(_03121_),
    .B1(_00360_),
    .Y(_05760_)
  );
  sg13g2_a21oi_1 _15704_ (
    .A1(_01029_),
    .A2(_05760_),
    .B1(_08487_),
    .Y(_05761_)
  );
  sg13g2_nor2_1 _15705_ (
    .A(_05759_),
    .B(_05761_),
    .Y(_05762_)
  );
  sg13g2_nor2_1 _15706_ (
    .A(_07171_),
    .B(_01064_),
    .Y(_05763_)
  );
  sg13g2_a21oi_1 _15707_ (
    .A1(_01507_),
    .A2(_00376_),
    .B1(_05575_),
    .Y(_05764_)
  );
  sg13g2_nor2_1 _15708_ (
    .A(_00678_),
    .B(_03709_),
    .Y(_05765_)
  );
  sg13g2_a22oi_1 _15709_ (
    .A1(_01472_),
    .A2(_00209_),
    .B1(_01627_),
    .B2(_05765_),
    .Y(_05766_)
  );
  sg13g2_nand3_1 _15710_ (
    .A(_05763_),
    .B(_05764_),
    .C(_05766_),
    .Y(_05768_)
  );
  sg13g2_nor2_1 _15711_ (
    .A(addr_i_2_),
    .B(_07038_),
    .Y(_05769_)
  );
  sg13g2_o21ai_1 _15712_ (
    .A1(_02204_),
    .A2(_05769_),
    .B1(addr_i_4_),
    .Y(_05770_)
  );
  sg13g2_nand3_1 _15713_ (
    .A(addr_i_3_),
    .B(_01331_),
    .C(_05770_),
    .Y(_05771_)
  );
  sg13g2_o21ai_1 _15714_ (
    .A1(addr_i_3_),
    .A2(_05768_),
    .B1(_05771_),
    .Y(_05772_)
  );
  sg13g2_nand2_1 _15715_ (
    .A(_02344_),
    .B(_02874_),
    .Y(_05773_)
  );
  sg13g2_a21oi_1 _15716_ (
    .A1(_05629_),
    .A2(_05773_),
    .B1(_00629_),
    .Y(_05774_)
  );
  sg13g2_o21ai_1 _15717_ (
    .A1(_00400_),
    .A2(_01402_),
    .B1(addr_i_3_),
    .Y(_05775_)
  );
  sg13g2_nand4_1 _15718_ (
    .A(_00276_),
    .B(_02167_),
    .C(_05698_),
    .D(_05775_),
    .Y(_05776_)
  );
  sg13g2_nand2_1 _15719_ (
    .A(addr_i_9_),
    .B(_05776_),
    .Y(_05777_)
  );
  sg13g2_o21ai_1 _15720_ (
    .A1(_02268_),
    .A2(_03455_),
    .B1(addr_i_3_),
    .Y(_05779_)
  );
  sg13g2_nand2_1 _15721_ (
    .A(addr_i_4_),
    .B(_00890_),
    .Y(_05780_)
  );
  sg13g2_a21oi_1 _15722_ (
    .A1(_06088_),
    .A2(_05780_),
    .B1(addr_i_3_),
    .Y(_05781_)
  );
  sg13g2_a21oi_1 _15723_ (
    .A1(addr_i_6_),
    .A2(_03323_),
    .B1(_05781_),
    .Y(_05782_)
  );
  sg13g2_a21oi_1 _15724_ (
    .A1(_05779_),
    .A2(_05782_),
    .B1(_01034_),
    .Y(_05783_)
  );
  sg13g2_a22oi_1 _15725_ (
    .A1(_05772_),
    .A2(_05774_),
    .B1(_05777_),
    .B2(_05783_),
    .Y(_05784_)
  );
  sg13g2_a21oi_1 _15726_ (
    .A1(_05754_),
    .A2(_05762_),
    .B1(_05784_),
    .Y(_05785_)
  );
  sg13g2_o21ai_1 _15727_ (
    .A1(addr_i_10_),
    .A2(_05785_),
    .B1(addr_i_11_),
    .Y(_05786_)
  );
  sg13g2_o21ai_1 _15728_ (
    .A1(_06298_),
    .A2(_01106_),
    .B1(_06364_),
    .Y(_05787_)
  );
  sg13g2_nand2b_1 _15729_ (
    .A_N(_00911_),
    .B(addr_i_4_),
    .Y(_05788_)
  );
  sg13g2_nand3_1 _15730_ (
    .A(addr_i_3_),
    .B(_05787_),
    .C(_05788_),
    .Y(_05790_)
  );
  sg13g2_nand2_1 _15731_ (
    .A(_00019_),
    .B(_01353_),
    .Y(_05791_)
  );
  sg13g2_a22oi_1 _15732_ (
    .A1(addr_i_4_),
    .A2(_05791_),
    .B1(_07193_),
    .B2(addr_i_3_),
    .Y(_05792_)
  );
  sg13g2_nor2_1 _15733_ (
    .A(_01011_),
    .B(_05792_),
    .Y(_05793_)
  );
  sg13g2_nor3_1 _15734_ (
    .A(addr_i_3_),
    .B(_03446_),
    .C(_01022_),
    .Y(_05794_)
  );
  sg13g2_o21ai_1 _15735_ (
    .A1(_00280_),
    .A2(_05794_),
    .B1(addr_i_2_),
    .Y(_05795_)
  );
  sg13g2_a21oi_1 _15736_ (
    .A1(_01943_),
    .A2(_03942_),
    .B1(_06519_),
    .Y(_05796_)
  );
  sg13g2_a21oi_1 _15737_ (
    .A1(_05795_),
    .A2(_05796_),
    .B1(_07591_),
    .Y(_05797_)
  );
  sg13g2_a21oi_1 _15738_ (
    .A1(_05790_),
    .A2(_05793_),
    .B1(_05797_),
    .Y(_05798_)
  );
  sg13g2_nand3_1 _15739_ (
    .A(addr_i_6_),
    .B(_04222_),
    .C(_00816_),
    .Y(_05799_)
  );
  sg13g2_a21oi_1 _15740_ (
    .A1(_00819_),
    .A2(_02750_),
    .B1(_01274_),
    .Y(_05801_)
  );
  sg13g2_nor2_1 _15741_ (
    .A(_02304_),
    .B(_05544_),
    .Y(_05802_)
  );
  sg13g2_nand2b_1 _15742_ (
    .A_N(_02178_),
    .B(_09475_),
    .Y(_05803_)
  );
  sg13g2_o21ai_1 _15743_ (
    .A1(_05802_),
    .A2(_05803_),
    .B1(addr_i_9_),
    .Y(_05804_)
  );
  sg13g2_xnor2_1 _15744_ (
    .A(addr_i_3_),
    .B(_01461_),
    .Y(_05805_)
  );
  sg13g2_nor2_1 _15745_ (
    .A(addr_i_5_),
    .B(_05805_),
    .Y(_05806_)
  );
  sg13g2_nor3_1 _15746_ (
    .A(_04661_),
    .B(_01746_),
    .C(_05806_),
    .Y(_05807_)
  );
  sg13g2_a22oi_1 _15747_ (
    .A1(_05799_),
    .A2(_05801_),
    .B1(_05804_),
    .B2(_05807_),
    .Y(_05808_)
  );
  sg13g2_o21ai_1 _15748_ (
    .A1(_01896_),
    .A2(_03188_),
    .B1(addr_i_4_),
    .Y(_05809_)
  );
  sg13g2_nor4_1 _15749_ (
    .A(_00547_),
    .B(_07967_),
    .C(_01659_),
    .D(_07270_),
    .Y(_05810_)
  );
  sg13g2_a22oi_1 _15750_ (
    .A1(_09473_),
    .A2(_05809_),
    .B1(_05810_),
    .B2(_01610_),
    .Y(_05812_)
  );
  sg13g2_nor2_1 _15751_ (
    .A(_08343_),
    .B(_09509_),
    .Y(_05813_)
  );
  sg13g2_a221oi_1 _15752_ (
    .A1(addr_i_4_),
    .A2(_07061_),
    .B1(_03413_),
    .B2(_07237_),
    .C1(_07712_),
    .Y(_05814_)
  );
  sg13g2_nor2_1 _15753_ (
    .A(addr_i_7_),
    .B(_01153_),
    .Y(_05815_)
  );
  sg13g2_a22oi_1 _15754_ (
    .A1(_01113_),
    .A2(_05815_),
    .B1(_01659_),
    .B2(addr_i_3_),
    .Y(_05816_)
  );
  sg13g2_a21oi_1 _15755_ (
    .A1(addr_i_3_),
    .A2(_05814_),
    .B1(_05816_),
    .Y(_05817_)
  );
  sg13g2_o21ai_1 _15756_ (
    .A1(_05813_),
    .A2(_05817_),
    .B1(addr_i_6_),
    .Y(_05818_)
  );
  sg13g2_nand2_1 _15757_ (
    .A(addr_i_3_),
    .B(_02241_),
    .Y(_05819_)
  );
  sg13g2_o21ai_1 _15758_ (
    .A1(_01153_),
    .A2(_01910_),
    .B1(_08741_),
    .Y(_05820_)
  );
  sg13g2_a21oi_1 _15759_ (
    .A1(_05819_),
    .A2(_05820_),
    .B1(_00505_),
    .Y(_05821_)
  );
  sg13g2_nand2_1 _15760_ (
    .A(_01384_),
    .B(_02218_),
    .Y(_05823_)
  );
  sg13g2_a22oi_1 _15761_ (
    .A1(_05302_),
    .A2(_05823_),
    .B1(_01041_),
    .B2(_00052_),
    .Y(_05824_)
  );
  sg13g2_a221oi_1 _15762_ (
    .A1(_03288_),
    .A2(_00650_),
    .B1(_01309_),
    .B2(_00534_),
    .C1(addr_i_7_),
    .Y(_05825_)
  );
  sg13g2_nor4_1 _15763_ (
    .A(_00213_),
    .B(_05821_),
    .C(_05824_),
    .D(_05825_),
    .Y(_05826_)
  );
  sg13g2_a221oi_1 _15764_ (
    .A1(_05798_),
    .A2(_05808_),
    .B1(_05812_),
    .B2(_05818_),
    .C1(_05826_),
    .Y(_05827_)
  );
  sg13g2_nor2_1 _15765_ (
    .A(addr_i_10_),
    .B(_05827_),
    .Y(_05828_)
  );
  sg13g2_o21ai_1 _15766_ (
    .A1(_01616_),
    .A2(_02742_),
    .B1(_04191_),
    .Y(_05829_)
  );
  sg13g2_a22oi_1 _15767_ (
    .A1(_03263_),
    .A2(_07679_),
    .B1(_01957_),
    .B2(addr_i_4_),
    .Y(_05830_)
  );
  sg13g2_a22oi_1 _15768_ (
    .A1(addr_i_4_),
    .A2(_05829_),
    .B1(_05830_),
    .B2(_01034_),
    .Y(_05831_)
  );
  sg13g2_a221oi_1 _15769_ (
    .A1(_01047_),
    .A2(_00226_),
    .B1(_02498_),
    .B2(_01888_),
    .C1(addr_i_3_),
    .Y(_05832_)
  );
  sg13g2_a221oi_1 _15770_ (
    .A1(_01047_),
    .A2(_02141_),
    .B1(_02498_),
    .B2(_08696_),
    .C1(_01067_),
    .Y(_05835_)
  );
  sg13g2_nor2_1 _15771_ (
    .A(_05832_),
    .B(_05835_),
    .Y(_05836_)
  );
  sg13g2_a22oi_1 _15772_ (
    .A1(_08951_),
    .A2(_03556_),
    .B1(_08056_),
    .B2(_00715_),
    .Y(_05837_)
  );
  sg13g2_a21oi_1 _15773_ (
    .A1(_01175_),
    .A2(_04093_),
    .B1(addr_i_4_),
    .Y(_05838_)
  );
  sg13g2_nor4_1 _15774_ (
    .A(_01494_),
    .B(_00494_),
    .C(_00885_),
    .D(_05838_),
    .Y(_05839_)
  );
  sg13g2_nor2_1 _15775_ (
    .A(_02459_),
    .B(_03132_),
    .Y(_05840_)
  );
  sg13g2_a21oi_1 _15776_ (
    .A1(addr_i_2_),
    .A2(_01047_),
    .B1(_05840_),
    .Y(_05841_)
  );
  sg13g2_nor3_1 _15777_ (
    .A(_01896_),
    .B(_02179_),
    .C(_04130_),
    .Y(_05842_)
  );
  sg13g2_a22oi_1 _15778_ (
    .A1(_06220_),
    .A2(_02498_),
    .B1(_05842_),
    .B2(_03073_),
    .Y(_05843_)
  );
  sg13g2_o21ai_1 _15779_ (
    .A1(addr_i_4_),
    .A2(_05841_),
    .B1(_05843_),
    .Y(_05844_)
  );
  sg13g2_nor4_1 _15780_ (
    .A(_05836_),
    .B(_05837_),
    .C(_05839_),
    .D(_05844_),
    .Y(_05846_)
  );
  sg13g2_nor2b_1 _15781_ (
    .A(_05831_),
    .B_N(_05846_),
    .Y(_05847_)
  );
  sg13g2_a22oi_1 _15782_ (
    .A1(addr_i_5_),
    .A2(_02505_),
    .B1(_02772_),
    .B2(_00060_),
    .Y(_05848_)
  );
  sg13g2_nor3_1 _15783_ (
    .A(addr_i_3_),
    .B(_04683_),
    .C(_00305_),
    .Y(_05849_)
  );
  sg13g2_a21oi_1 _15784_ (
    .A1(_09205_),
    .A2(_00138_),
    .B1(addr_i_4_),
    .Y(_05850_)
  );
  sg13g2_nor2_1 _15785_ (
    .A(addr_i_7_),
    .B(_05850_),
    .Y(_05851_)
  );
  sg13g2_o21ai_1 _15786_ (
    .A1(_05848_),
    .A2(_05849_),
    .B1(_05851_),
    .Y(_05852_)
  );
  sg13g2_nand2_1 _15787_ (
    .A(_08254_),
    .B(_08951_),
    .Y(_05853_)
  );
  sg13g2_a21oi_1 _15788_ (
    .A1(_00573_),
    .A2(_03927_),
    .B1(addr_i_3_),
    .Y(_05854_)
  );
  sg13g2_nand2_1 _15789_ (
    .A(addr_i_7_),
    .B(_00118_),
    .Y(_05855_)
  );
  sg13g2_a22oi_1 _15790_ (
    .A1(addr_i_2_),
    .A2(_05853_),
    .B1(_05854_),
    .B2(_05855_),
    .Y(_05857_)
  );
  sg13g2_nor2_1 _15791_ (
    .A(addr_i_8_),
    .B(_05857_),
    .Y(_05858_)
  );
  sg13g2_o21ai_1 _15792_ (
    .A1(_01910_),
    .A2(_02322_),
    .B1(addr_i_3_),
    .Y(_05859_)
  );
  sg13g2_nand2_1 _15793_ (
    .A(_01230_),
    .B(_05859_),
    .Y(_05860_)
  );
  sg13g2_o21ai_1 _15794_ (
    .A1(_00377_),
    .A2(_00234_),
    .B1(_00159_),
    .Y(_05861_)
  );
  sg13g2_a21oi_1 _15795_ (
    .A1(_03853_),
    .A2(_00808_),
    .B1(_00112_),
    .Y(_05862_)
  );
  sg13g2_nand2_1 _15796_ (
    .A(_05861_),
    .B(_05862_),
    .Y(_05863_)
  );
  sg13g2_nand2_1 _15797_ (
    .A(_06088_),
    .B(_05243_),
    .Y(_05864_)
  );
  sg13g2_nor2_1 _15798_ (
    .A(_02404_),
    .B(_01031_),
    .Y(_05865_)
  );
  sg13g2_nor3_1 _15799_ (
    .A(addr_i_3_),
    .B(_07359_),
    .C(_01660_),
    .Y(_05866_)
  );
  sg13g2_a22oi_1 _15800_ (
    .A1(_05864_),
    .A2(_05865_),
    .B1(_05866_),
    .B2(_05822_),
    .Y(_05868_)
  );
  sg13g2_a22oi_1 _15801_ (
    .A1(_02257_),
    .A2(_05860_),
    .B1(_05863_),
    .B2(_05868_),
    .Y(_05869_)
  );
  sg13g2_a22oi_1 _15802_ (
    .A1(_05852_),
    .A2(_05858_),
    .B1(_05869_),
    .B2(_00925_),
    .Y(_05870_)
  );
  sg13g2_or4_1 _15803_ (
    .A(addr_i_11_),
    .B(_05828_),
    .C(_05847_),
    .D(_05870_),
    .X(_05871_)
  );
  sg13g2_o21ai_1 _15804_ (
    .A1(_05743_),
    .A2(_05786_),
    .B1(_05871_),
    .Y(_05872_)
  );
  sg13g2_mux2_1 _15805_ (
    .A0(_05703_),
    .A1(_05872_),
    .S(_02251_),
    .X(data_o_25_)
  );
  sg13g2_nand2_1 _15806_ (
    .A(_00150_),
    .B(_09478_),
    .Y(_05873_)
  );
  sg13g2_a221oi_1 _15807_ (
    .A1(addr_i_6_),
    .A2(_05873_),
    .B1(_02585_),
    .B2(addr_i_3_),
    .C1(_00084_),
    .Y(_05874_)
  );
  sg13g2_a22oi_1 _15808_ (
    .A1(_03431_),
    .A2(_00999_),
    .B1(_00824_),
    .B2(addr_i_4_),
    .Y(_05875_)
  );
  sg13g2_o21ai_1 _15809_ (
    .A1(_05874_),
    .A2(_05875_),
    .B1(addr_i_7_),
    .Y(_05876_)
  );
  sg13g2_a21oi_1 _15810_ (
    .A1(_03431_),
    .A2(_00820_),
    .B1(addr_i_4_),
    .Y(_05878_)
  );
  sg13g2_nor2_1 _15811_ (
    .A(_00390_),
    .B(_05878_),
    .Y(_05879_)
  );
  sg13g2_a22oi_1 _15812_ (
    .A1(_00617_),
    .A2(_07911_),
    .B1(_01481_),
    .B2(_04442_),
    .Y(_05880_)
  );
  sg13g2_a22oi_1 _15813_ (
    .A1(_03182_),
    .A2(_05879_),
    .B1(_05880_),
    .B2(addr_i_8_),
    .Y(_05881_)
  );
  sg13g2_o21ai_1 _15814_ (
    .A1(addr_i_2_),
    .A2(_01262_),
    .B1(_00626_),
    .Y(_05882_)
  );
  sg13g2_nor2_1 _15815_ (
    .A(_07326_),
    .B(_00547_),
    .Y(_05883_)
  );
  sg13g2_a21oi_1 _15816_ (
    .A1(addr_i_5_),
    .A2(_03358_),
    .B1(_03930_),
    .Y(_05884_)
  );
  sg13g2_nor2_1 _15817_ (
    .A(_05883_),
    .B(_05884_),
    .Y(_05885_)
  );
  sg13g2_nand2_1 _15818_ (
    .A(_05882_),
    .B(_05885_),
    .Y(_05886_)
  );
  sg13g2_o21ai_1 _15819_ (
    .A1(_02265_),
    .A2(_09499_),
    .B1(_01336_),
    .Y(_05887_)
  );
  sg13g2_a22oi_1 _15820_ (
    .A1(addr_i_4_),
    .A2(_00476_),
    .B1(_00632_),
    .B2(_01169_),
    .Y(_05889_)
  );
  sg13g2_o21ai_1 _15821_ (
    .A1(addr_i_5_),
    .A2(_01326_),
    .B1(_05889_),
    .Y(_05890_)
  );
  sg13g2_nand4_1 _15822_ (
    .A(addr_i_8_),
    .B(_00658_),
    .C(_05887_),
    .D(_05890_),
    .Y(_05891_)
  );
  sg13g2_a21oi_1 _15823_ (
    .A1(addr_i_4_),
    .A2(_05886_),
    .B1(_05891_),
    .Y(_05892_)
  );
  sg13g2_a22oi_1 _15824_ (
    .A1(_05876_),
    .A2(_05881_),
    .B1(_05892_),
    .B2(_00109_),
    .Y(_05893_)
  );
  sg13g2_a21oi_1 _15825_ (
    .A1(_05888_),
    .A2(_06895_),
    .B1(_02297_),
    .Y(_05894_)
  );
  sg13g2_nor2_1 _15826_ (
    .A(addr_i_4_),
    .B(_05107_),
    .Y(_05895_)
  );
  sg13g2_a22oi_1 _15827_ (
    .A1(addr_i_4_),
    .A2(_02781_),
    .B1(_05895_),
    .B2(_00067_),
    .Y(_05896_)
  );
  sg13g2_a22oi_1 _15828_ (
    .A1(addr_i_8_),
    .A2(_00128_),
    .B1(_05894_),
    .B2(_05896_),
    .Y(_05897_)
  );
  sg13g2_nand2b_1 _15829_ (
    .A_N(addr_i_8_),
    .B(addr_i_4_),
    .Y(_05898_)
  );
  sg13g2_nand3_1 _15830_ (
    .A(addr_i_5_),
    .B(_01914_),
    .C(_05898_),
    .Y(_05900_)
  );
  sg13g2_o21ai_1 _15831_ (
    .A1(addr_i_5_),
    .A2(_05898_),
    .B1(_05900_),
    .Y(_05901_)
  );
  sg13g2_nand2_1 _15832_ (
    .A(addr_i_2_),
    .B(addr_i_8_),
    .Y(_05902_)
  );
  sg13g2_nand2_1 _15833_ (
    .A(addr_i_4_),
    .B(_06331_),
    .Y(_05903_)
  );
  sg13g2_a21oi_1 _15834_ (
    .A1(_05902_),
    .A2(_05903_),
    .B1(_02777_),
    .Y(_05904_)
  );
  sg13g2_a21o_1 _15835_ (
    .A1(_08598_),
    .A2(_02781_),
    .B1(_05904_),
    .X(_05905_)
  );
  sg13g2_a22oi_1 _15836_ (
    .A1(addr_i_2_),
    .A2(_05901_),
    .B1(_05905_),
    .B2(addr_i_3_),
    .Y(_05906_)
  );
  sg13g2_a21oi_1 _15837_ (
    .A1(addr_i_3_),
    .A2(_05897_),
    .B1(_05906_),
    .Y(_05907_)
  );
  sg13g2_o21ai_1 _15838_ (
    .A1(_04952_),
    .A2(_05907_),
    .B1(addr_i_7_),
    .Y(_05908_)
  );
  sg13g2_a21oi_1 _15839_ (
    .A1(addr_i_6_),
    .A2(_01208_),
    .B1(_01308_),
    .Y(_05909_)
  );
  sg13g2_nor2_1 _15840_ (
    .A(addr_i_4_),
    .B(_05909_),
    .Y(_05911_)
  );
  sg13g2_nand2_1 _15841_ (
    .A(_02815_),
    .B(_01060_),
    .Y(_05912_)
  );
  sg13g2_a22oi_1 _15842_ (
    .A1(_00067_),
    .A2(_05912_),
    .B1(_01863_),
    .B2(_00659_),
    .Y(_05913_)
  );
  sg13g2_a22oi_1 _15843_ (
    .A1(_03521_),
    .A2(_05911_),
    .B1(_05913_),
    .B2(addr_i_8_),
    .Y(_05914_)
  );
  sg13g2_a21oi_1 _15844_ (
    .A1(_09510_),
    .A2(_05756_),
    .B1(addr_i_3_),
    .Y(_05915_)
  );
  sg13g2_o21ai_1 _15845_ (
    .A1(_04121_),
    .A2(_05915_),
    .B1(addr_i_4_),
    .Y(_05916_)
  );
  sg13g2_nand3_1 _15846_ (
    .A(_01104_),
    .B(_01257_),
    .C(_00157_),
    .Y(_05917_)
  );
  sg13g2_a21oi_1 _15847_ (
    .A1(_05916_),
    .A2(_05917_),
    .B1(_00782_),
    .Y(_05918_)
  );
  sg13g2_or3_1 _15848_ (
    .A(addr_i_7_),
    .B(_05914_),
    .C(_05918_),
    .X(_05919_)
  );
  sg13g2_a21oi_1 _15849_ (
    .A1(_05908_),
    .A2(_05919_),
    .B1(_01211_),
    .Y(_05920_)
  );
  sg13g2_nand2_1 _15850_ (
    .A(_00010_),
    .B(_01215_),
    .Y(_05922_)
  );
  sg13g2_a21oi_1 _15851_ (
    .A1(_00025_),
    .A2(_01221_),
    .B1(addr_i_2_),
    .Y(_05923_)
  );
  sg13g2_o21ai_1 _15852_ (
    .A1(_00297_),
    .A2(_05923_),
    .B1(addr_i_4_),
    .Y(_05924_)
  );
  sg13g2_o21ai_1 _15853_ (
    .A1(_09127_),
    .A2(_02632_),
    .B1(addr_i_2_),
    .Y(_05925_)
  );
  sg13g2_nand3_1 _15854_ (
    .A(_05922_),
    .B(_05924_),
    .C(_05925_),
    .Y(_05926_)
  );
  sg13g2_nand2_1 _15855_ (
    .A(_06364_),
    .B(_04429_),
    .Y(_05927_)
  );
  sg13g2_nor2_1 _15856_ (
    .A(_02623_),
    .B(_02634_),
    .Y(_05928_)
  );
  sg13g2_a21oi_1 _15857_ (
    .A1(addr_i_5_),
    .A2(_05927_),
    .B1(_05928_),
    .Y(_05929_)
  );
  sg13g2_o21ai_1 _15858_ (
    .A1(addr_i_3_),
    .A2(_05929_),
    .B1(_03420_),
    .Y(_05930_)
  );
  sg13g2_a21oi_1 _15859_ (
    .A1(_00650_),
    .A2(_05689_),
    .B1(_03743_),
    .Y(_05931_)
  );
  sg13g2_o21ai_1 _15860_ (
    .A1(_02424_),
    .A2(_05931_),
    .B1(_00778_),
    .Y(_05933_)
  );
  sg13g2_nand3_1 _15861_ (
    .A(_01559_),
    .B(_01740_),
    .C(_05933_),
    .Y(_05934_)
  );
  sg13g2_a221oi_1 _15862_ (
    .A1(addr_i_3_),
    .A2(_05926_),
    .B1(_05930_),
    .B2(addr_i_2_),
    .C1(_05934_),
    .Y(_05935_)
  );
  sg13g2_nand2_1 _15863_ (
    .A(addr_i_6_),
    .B(_02471_),
    .Y(_05936_)
  );
  sg13g2_a22oi_1 _15864_ (
    .A1(_09491_),
    .A2(_05936_),
    .B1(_00334_),
    .B2(_01231_),
    .Y(_05937_)
  );
  sg13g2_nand2_1 _15865_ (
    .A(_00258_),
    .B(_01223_),
    .Y(_05938_)
  );
  sg13g2_o21ai_1 _15866_ (
    .A1(addr_i_4_),
    .A2(_05937_),
    .B1(_05938_),
    .Y(_05939_)
  );
  sg13g2_a21oi_1 _15867_ (
    .A1(addr_i_2_),
    .A2(_02874_),
    .B1(_00132_),
    .Y(_05940_)
  );
  sg13g2_o21ai_1 _15868_ (
    .A1(addr_i_3_),
    .A2(_05940_),
    .B1(_01180_),
    .Y(_05941_)
  );
  sg13g2_a21oi_1 _15869_ (
    .A1(_06088_),
    .A2(_01420_),
    .B1(_00999_),
    .Y(_05942_)
  );
  sg13g2_o21ai_1 _15870_ (
    .A1(addr_i_7_),
    .A2(_05942_),
    .B1(addr_i_8_),
    .Y(_05945_)
  );
  sg13g2_a22oi_1 _15871_ (
    .A1(_00123_),
    .A2(_05939_),
    .B1(_05941_),
    .B2(_05945_),
    .Y(_05946_)
  );
  sg13g2_or3_1 _15872_ (
    .A(addr_i_9_),
    .B(_05935_),
    .C(_05946_),
    .X(_05947_)
  );
  sg13g2_a21oi_1 _15873_ (
    .A1(_01301_),
    .A2(_03457_),
    .B1(_00967_),
    .Y(_05948_)
  );
  sg13g2_o21ai_1 _15874_ (
    .A1(_00119_),
    .A2(_05948_),
    .B1(_00146_),
    .Y(_05949_)
  );
  sg13g2_a21oi_1 _15875_ (
    .A1(_08431_),
    .A2(_00417_),
    .B1(addr_i_3_),
    .Y(_05950_)
  );
  sg13g2_nor2_1 _15876_ (
    .A(addr_i_7_),
    .B(_05950_),
    .Y(_05951_)
  );
  sg13g2_o21ai_1 _15877_ (
    .A1(_02287_),
    .A2(_00412_),
    .B1(_01224_),
    .Y(_05952_)
  );
  sg13g2_nand2_1 _15878_ (
    .A(addr_i_7_),
    .B(_02167_),
    .Y(_05953_)
  );
  sg13g2_a21oi_1 _15879_ (
    .A1(addr_i_4_),
    .A2(_02858_),
    .B1(_01015_),
    .Y(_05954_)
  );
  sg13g2_nor2_1 _15880_ (
    .A(_02271_),
    .B(_05954_),
    .Y(_05956_)
  );
  sg13g2_a22oi_1 _15881_ (
    .A1(_01935_),
    .A2(_05952_),
    .B1(_05953_),
    .B2(_05956_),
    .Y(_05957_)
  );
  sg13g2_a22oi_1 _15882_ (
    .A1(_05949_),
    .A2(_05951_),
    .B1(_05957_),
    .B2(_01151_),
    .Y(_05958_)
  );
  sg13g2_nand2_1 _15883_ (
    .A(addr_i_4_),
    .B(_00282_),
    .Y(_05959_)
  );
  sg13g2_a21oi_1 _15884_ (
    .A1(addr_i_4_),
    .A2(_00327_),
    .B1(_07658_),
    .Y(_05960_)
  );
  sg13g2_nand2_1 _15885_ (
    .A(_00200_),
    .B(_05960_),
    .Y(_05961_)
  );
  sg13g2_a21oi_1 _15886_ (
    .A1(_05959_),
    .A2(_05961_),
    .B1(addr_i_3_),
    .Y(_05962_)
  );
  sg13g2_a221oi_1 _15887_ (
    .A1(_07547_),
    .A2(_00770_),
    .B1(_02166_),
    .B2(addr_i_3_),
    .C1(_05962_),
    .Y(_05963_)
  );
  sg13g2_nand2b_1 _15888_ (
    .A_N(_02943_),
    .B(_01674_),
    .Y(_05964_)
  );
  sg13g2_o21ai_1 _15889_ (
    .A1(addr_i_4_),
    .A2(_01459_),
    .B1(addr_i_3_),
    .Y(_05965_)
  );
  sg13g2_nand3_1 _15890_ (
    .A(_07625_),
    .B(_02002_),
    .C(_05965_),
    .Y(_05967_)
  );
  sg13g2_a221oi_1 _15891_ (
    .A1(_09138_),
    .A2(_05964_),
    .B1(_05967_),
    .B2(_01320_),
    .C1(addr_i_8_),
    .Y(_05968_)
  );
  sg13g2_o21ai_1 _15892_ (
    .A1(addr_i_7_),
    .A2(_05963_),
    .B1(_05968_),
    .Y(_05969_)
  );
  sg13g2_nand3b_1 _15893_ (
    .A_N(_05958_),
    .B(addr_i_9_),
    .C(_05969_),
    .Y(_05970_)
  );
  sg13g2_a21oi_1 _15894_ (
    .A1(_05947_),
    .A2(_05970_),
    .B1(addr_i_10_),
    .Y(_05971_)
  );
  sg13g2_nor4_1 _15895_ (
    .A(addr_i_11_),
    .B(_05893_),
    .C(_05920_),
    .D(_05971_),
    .Y(_05972_)
  );
  sg13g2_inv_1 _15896_ (
    .A(_00667_),
    .Y(_05973_)
  );
  sg13g2_a21oi_1 _15897_ (
    .A1(_00771_),
    .A2(_05973_),
    .B1(_00403_),
    .Y(_05974_)
  );
  sg13g2_a21oi_1 _15898_ (
    .A1(addr_i_7_),
    .A2(_05974_),
    .B1(_05833_),
    .Y(_05975_)
  );
  sg13g2_o21ai_1 _15899_ (
    .A1(_02040_),
    .A2(_05975_),
    .B1(addr_i_11_),
    .Y(_05976_)
  );
  sg13g2_a21o_1 _15900_ (
    .A1(_00172_),
    .A2(_03238_),
    .B1(_00201_),
    .X(_05978_)
  );
  sg13g2_o21ai_1 _15901_ (
    .A1(_03032_),
    .A2(_00266_),
    .B1(addr_i_2_),
    .Y(_05979_)
  );
  sg13g2_nand2_1 _15902_ (
    .A(_00779_),
    .B(_05979_),
    .Y(_05980_)
  );
  sg13g2_inv_1 _15903_ (
    .A(_02850_),
    .Y(_05981_)
  );
  sg13g2_a22oi_1 _15904_ (
    .A1(_00047_),
    .A2(_05981_),
    .B1(_02801_),
    .B2(_07370_),
    .Y(_05982_)
  );
  sg13g2_nor2_1 _15905_ (
    .A(_01481_),
    .B(_05982_),
    .Y(_05983_)
  );
  sg13g2_a22oi_1 _15906_ (
    .A1(_00172_),
    .A2(_05980_),
    .B1(_05983_),
    .B2(_06706_),
    .Y(_05984_)
  );
  sg13g2_nand2_1 _15907_ (
    .A(_00716_),
    .B(_00368_),
    .Y(_05985_)
  );
  sg13g2_a21oi_1 _15908_ (
    .A1(addr_i_6_),
    .A2(_01808_),
    .B1(addr_i_3_),
    .Y(_05986_)
  );
  sg13g2_a221oi_1 _15909_ (
    .A1(_09105_),
    .A2(_01500_),
    .B1(_05985_),
    .B2(addr_i_3_),
    .C1(_05986_),
    .Y(_05987_)
  );
  sg13g2_nand2_1 _15910_ (
    .A(_00150_),
    .B(_01265_),
    .Y(_05989_)
  );
  sg13g2_a21oi_1 _15911_ (
    .A1(_01257_),
    .A2(_03559_),
    .B1(addr_i_4_),
    .Y(_05990_)
  );
  sg13g2_a22oi_1 _15912_ (
    .A1(addr_i_3_),
    .A2(_05989_),
    .B1(_05990_),
    .B2(_01846_),
    .Y(_05991_)
  );
  sg13g2_nand2b_1 _15913_ (
    .A_N(_05991_),
    .B(_00610_),
    .Y(_05992_)
  );
  sg13g2_o21ai_1 _15914_ (
    .A1(_01082_),
    .A2(_05987_),
    .B1(_05992_),
    .Y(_05993_)
  );
  sg13g2_nor3_1 _15915_ (
    .A(addr_i_9_),
    .B(_05984_),
    .C(_05993_),
    .Y(_05994_)
  );
  sg13g2_a22oi_1 _15916_ (
    .A1(addr_i_9_),
    .A2(_05978_),
    .B1(_05994_),
    .B2(addr_i_10_),
    .Y(_05995_)
  );
  sg13g2_o21ai_1 _15917_ (
    .A1(_05976_),
    .A2(_05995_),
    .B1(addr_i_12_),
    .Y(_05996_)
  );
  sg13g2_a21oi_1 _15918_ (
    .A1(_03540_),
    .A2(_00442_),
    .B1(_02123_),
    .Y(_05997_)
  );
  sg13g2_o21ai_1 _15919_ (
    .A1(_05280_),
    .A2(_01747_),
    .B1(addr_i_4_),
    .Y(_05998_)
  );
  sg13g2_o21ai_1 _15920_ (
    .A1(addr_i_5_),
    .A2(_05997_),
    .B1(_05998_),
    .Y(_06000_)
  );
  sg13g2_o21ai_1 _15921_ (
    .A1(_01277_),
    .A2(_01571_),
    .B1(addr_i_4_),
    .Y(_06001_)
  );
  sg13g2_nand3_1 _15922_ (
    .A(_01212_),
    .B(_00155_),
    .C(_01571_),
    .Y(_06002_)
  );
  sg13g2_o21ai_1 _15923_ (
    .A1(_02976_),
    .A2(_03589_),
    .B1(addr_i_6_),
    .Y(_06003_)
  );
  sg13g2_nand3_1 _15924_ (
    .A(_06001_),
    .B(_06002_),
    .C(_06003_),
    .Y(_06004_)
  );
  sg13g2_a22oi_1 _15925_ (
    .A1(_00388_),
    .A2(_06000_),
    .B1(_06004_),
    .B2(addr_i_8_),
    .Y(_06005_)
  );
  sg13g2_a21o_1 _15926_ (
    .A1(addr_i_3_),
    .A2(_04613_),
    .B1(_04681_),
    .X(_06006_)
  );
  sg13g2_a21o_1 _15927_ (
    .A1(_00676_),
    .A2(_07492_),
    .B1(_01654_),
    .X(_06007_)
  );
  sg13g2_o21ai_1 _15928_ (
    .A1(_03908_),
    .A2(_03106_),
    .B1(_04450_),
    .Y(_06008_)
  );
  sg13g2_a21oi_1 _15929_ (
    .A1(_01422_),
    .A2(_06008_),
    .B1(addr_i_5_),
    .Y(_06009_)
  );
  sg13g2_o21ai_1 _15930_ (
    .A1(addr_i_2_),
    .A2(_00578_),
    .B1(_05811_),
    .Y(_06011_)
  );
  sg13g2_a22oi_1 _15931_ (
    .A1(addr_i_2_),
    .A2(_06007_),
    .B1(_06009_),
    .B2(_06011_),
    .Y(_06012_)
  );
  sg13g2_a22oi_1 _15932_ (
    .A1(addr_i_7_),
    .A2(_06006_),
    .B1(_06012_),
    .B2(_05266_),
    .Y(_06013_)
  );
  sg13g2_nor2_1 _15933_ (
    .A(_01043_),
    .B(_06013_),
    .Y(_06014_)
  );
  sg13g2_o21ai_1 _15934_ (
    .A1(_06005_),
    .A2(_06014_),
    .B1(addr_i_9_),
    .Y(_06015_)
  );
  sg13g2_nor2_1 _15935_ (
    .A(_09371_),
    .B(_06320_),
    .Y(_06016_)
  );
  sg13g2_nand2_1 _15936_ (
    .A(addr_i_8_),
    .B(addr_i_6_),
    .Y(_06017_)
  );
  sg13g2_nor3_1 _15937_ (
    .A(addr_i_2_),
    .B(_01920_),
    .C(_01936_),
    .Y(_06018_)
  );
  sg13g2_a22oi_1 _15938_ (
    .A1(addr_i_2_),
    .A2(_06017_),
    .B1(_06018_),
    .B2(_06143_),
    .Y(_06019_)
  );
  sg13g2_o21ai_1 _15939_ (
    .A1(_06016_),
    .A2(_06019_),
    .B1(addr_i_3_),
    .Y(_06020_)
  );
  sg13g2_a21oi_1 _15940_ (
    .A1(_00586_),
    .A2(_01928_),
    .B1(addr_i_5_),
    .Y(_06022_)
  );
  sg13g2_a21oi_1 _15941_ (
    .A1(_06342_),
    .A2(_02462_),
    .B1(_06022_),
    .Y(_06023_)
  );
  sg13g2_a21o_1 _15942_ (
    .A1(_06020_),
    .A2(_06023_),
    .B1(addr_i_4_),
    .X(_06024_)
  );
  sg13g2_o21ai_1 _15943_ (
    .A1(addr_i_3_),
    .A2(_05955_),
    .B1(_02218_),
    .Y(_06025_)
  );
  sg13g2_nand2_1 _15944_ (
    .A(addr_i_2_),
    .B(_01920_),
    .Y(_06026_)
  );
  sg13g2_o21ai_1 _15945_ (
    .A1(_00819_),
    .A2(_06026_),
    .B1(addr_i_4_),
    .Y(_06027_)
  );
  sg13g2_a21oi_1 _15946_ (
    .A1(_01175_),
    .A2(_01843_),
    .B1(addr_i_8_),
    .Y(_06028_)
  );
  sg13g2_a22oi_1 _15947_ (
    .A1(_00448_),
    .A2(_06025_),
    .B1(_06027_),
    .B2(_06028_),
    .Y(_06029_)
  );
  sg13g2_a22oi_1 _15948_ (
    .A1(_00223_),
    .A2(_06021_),
    .B1(_06029_),
    .B2(_00351_),
    .Y(_06030_)
  );
  sg13g2_nand2_1 _15949_ (
    .A(_00990_),
    .B(_07458_),
    .Y(_06031_)
  );
  sg13g2_nor2_1 _15950_ (
    .A(_08156_),
    .B(_00495_),
    .Y(_06033_)
  );
  sg13g2_o21ai_1 _15951_ (
    .A1(_03170_),
    .A2(_06033_),
    .B1(_05402_),
    .Y(_06034_)
  );
  sg13g2_a21oi_1 _15952_ (
    .A1(_06031_),
    .A2(_06034_),
    .B1(_00112_),
    .Y(_06035_)
  );
  sg13g2_o21ai_1 _15953_ (
    .A1(_05524_),
    .A2(_06198_),
    .B1(_06143_),
    .Y(_06036_)
  );
  sg13g2_o21ai_1 _15954_ (
    .A1(addr_i_8_),
    .A2(_07658_),
    .B1(_07757_),
    .Y(_06037_)
  );
  sg13g2_a21oi_1 _15955_ (
    .A1(_05902_),
    .A2(_01033_),
    .B1(addr_i_3_),
    .Y(_06038_)
  );
  sg13g2_nand4_1 _15956_ (
    .A(_06026_),
    .B(_06036_),
    .C(_06037_),
    .D(_06038_),
    .Y(_06039_)
  );
  sg13g2_nand4_1 _15957_ (
    .A(addr_i_3_),
    .B(_01548_),
    .C(_00079_),
    .D(_00702_),
    .Y(_06040_)
  );
  sg13g2_nand3_1 _15958_ (
    .A(_06619_),
    .B(_06039_),
    .C(_06040_),
    .Y(_06041_)
  );
  sg13g2_nor2_1 _15959_ (
    .A(_06035_),
    .B(_06041_),
    .Y(_06042_)
  );
  sg13g2_a22oi_1 _15960_ (
    .A1(_06024_),
    .A2(_06030_),
    .B1(_06042_),
    .B2(addr_i_9_),
    .Y(_06044_)
  );
  sg13g2_nor2_1 _15961_ (
    .A(addr_i_10_),
    .B(_06044_),
    .Y(_06045_)
  );
  sg13g2_o21ai_1 _15962_ (
    .A1(_01582_),
    .A2(_02330_),
    .B1(addr_i_5_),
    .Y(_06046_)
  );
  sg13g2_a22oi_1 _15963_ (
    .A1(_07824_),
    .A2(_01813_),
    .B1(_00206_),
    .B2(addr_i_7_),
    .Y(_06047_)
  );
  sg13g2_nand2_1 _15964_ (
    .A(_00239_),
    .B(_01635_),
    .Y(_06048_)
  );
  sg13g2_nand3_1 _15965_ (
    .A(_06046_),
    .B(_06047_),
    .C(_06048_),
    .Y(_06049_)
  );
  sg13g2_o21ai_1 _15966_ (
    .A1(_07911_),
    .A2(_00544_),
    .B1(_00168_),
    .Y(_06050_)
  );
  sg13g2_or2_1 _15967_ (
    .A(_01536_),
    .B(_06050_),
    .X(_06051_)
  );
  sg13g2_nand2_1 _15968_ (
    .A(addr_i_3_),
    .B(_04186_),
    .Y(_06052_)
  );
  sg13g2_nand3_1 _15969_ (
    .A(_00529_),
    .B(_09476_),
    .C(_06052_),
    .Y(_06053_)
  );
  sg13g2_nand4_1 _15970_ (
    .A(addr_i_8_),
    .B(_06049_),
    .C(_06051_),
    .D(_06053_),
    .Y(_06056_)
  );
  sg13g2_a21oi_1 _15971_ (
    .A1(_00747_),
    .A2(_06508_),
    .B1(_00324_),
    .Y(_06057_)
  );
  sg13g2_nand2_1 _15972_ (
    .A(_00930_),
    .B(_01244_),
    .Y(_06058_)
  );
  sg13g2_o21ai_1 _15973_ (
    .A1(_00716_),
    .A2(_01747_),
    .B1(_06058_),
    .Y(_06059_)
  );
  sg13g2_o21ai_1 _15974_ (
    .A1(_00844_),
    .A2(_03358_),
    .B1(_01005_),
    .Y(_06060_)
  );
  sg13g2_a22oi_1 _15975_ (
    .A1(addr_i_2_),
    .A2(_06059_),
    .B1(_06060_),
    .B2(addr_i_6_),
    .Y(_06061_)
  );
  sg13g2_a221oi_1 _15976_ (
    .A1(_00861_),
    .A2(_00972_),
    .B1(_00727_),
    .B2(_02404_),
    .C1(_02685_),
    .Y(_06062_)
  );
  sg13g2_nor2_1 _15977_ (
    .A(_00825_),
    .B(_06062_),
    .Y(_06063_)
  );
  sg13g2_nor4_1 _15978_ (
    .A(addr_i_8_),
    .B(_06057_),
    .C(_06061_),
    .D(_06063_),
    .Y(_06064_)
  );
  sg13g2_nor2_1 _15979_ (
    .A(_03073_),
    .B(_06064_),
    .Y(_06065_)
  );
  sg13g2_o21ai_1 _15980_ (
    .A1(addr_i_4_),
    .A2(_00014_),
    .B1(addr_i_3_),
    .Y(_06067_)
  );
  sg13g2_o21ai_1 _15981_ (
    .A1(addr_i_2_),
    .A2(_03695_),
    .B1(_06067_),
    .Y(_06068_)
  );
  sg13g2_a221oi_1 _15982_ (
    .A1(_00319_),
    .A2(_02626_),
    .B1(_03046_),
    .B2(_04539_),
    .C1(addr_i_7_),
    .Y(_06069_)
  );
  sg13g2_nand2_1 _15983_ (
    .A(_00044_),
    .B(_03490_),
    .Y(_06070_)
  );
  sg13g2_a21oi_1 _15984_ (
    .A1(addr_i_3_),
    .A2(_06070_),
    .B1(_00304_),
    .Y(_06071_)
  );
  sg13g2_nand2b_1 _15985_ (
    .A_N(_06071_),
    .B(addr_i_5_),
    .Y(_06072_)
  );
  sg13g2_a21oi_1 _15986_ (
    .A1(_03089_),
    .A2(_05334_),
    .B1(_00505_),
    .Y(_06073_)
  );
  sg13g2_a221oi_1 _15987_ (
    .A1(_00168_),
    .A2(_06068_),
    .B1(_06069_),
    .B2(_06072_),
    .C1(_06073_),
    .Y(_06074_)
  );
  sg13g2_a21oi_1 _15988_ (
    .A1(_01175_),
    .A2(_00358_),
    .B1(_05302_),
    .Y(_06075_)
  );
  sg13g2_o21ai_1 _15989_ (
    .A1(_02733_),
    .A2(_03045_),
    .B1(_01353_),
    .Y(_06076_)
  );
  sg13g2_a22oi_1 _15990_ (
    .A1(_00726_),
    .A2(_02585_),
    .B1(_06075_),
    .B2(_06076_),
    .Y(_06078_)
  );
  sg13g2_o21ai_1 _15991_ (
    .A1(addr_i_2_),
    .A2(_03695_),
    .B1(_00993_),
    .Y(_06079_)
  );
  sg13g2_a221oi_1 _15992_ (
    .A1(_06099_),
    .A2(_00224_),
    .B1(_05634_),
    .B2(_02746_),
    .C1(_00780_),
    .Y(_06080_)
  );
  sg13g2_a21oi_1 _15993_ (
    .A1(_06079_),
    .A2(_06080_),
    .B1(_00108_),
    .Y(_06081_)
  );
  sg13g2_o21ai_1 _15994_ (
    .A1(_00860_),
    .A2(_06078_),
    .B1(_06081_),
    .Y(_06082_)
  );
  sg13g2_a21oi_1 _15995_ (
    .A1(addr_i_8_),
    .A2(_06074_),
    .B1(_06082_),
    .Y(_06083_)
  );
  sg13g2_nand2b_1 _15996_ (
    .A_N(_06083_),
    .B(addr_i_11_),
    .Y(_06084_)
  );
  sg13g2_a221oi_1 _15997_ (
    .A1(_06015_),
    .A2(_06045_),
    .B1(_06056_),
    .B2(_06065_),
    .C1(_06084_),
    .Y(_06085_)
  );
  sg13g2_a21oi_1 _15998_ (
    .A1(_00736_),
    .A2(_02001_),
    .B1(addr_i_4_),
    .Y(_06086_)
  );
  sg13g2_a21oi_1 _15999_ (
    .A1(_09161_),
    .A2(_00039_),
    .B1(addr_i_3_),
    .Y(_06087_)
  );
  sg13g2_a22oi_1 _16000_ (
    .A1(addr_i_3_),
    .A2(_03932_),
    .B1(_06086_),
    .B2(_06087_),
    .Y(_06089_)
  );
  sg13g2_nor2_1 _16001_ (
    .A(addr_i_7_),
    .B(_06089_),
    .Y(_06090_)
  );
  sg13g2_a22oi_1 _16002_ (
    .A1(_03431_),
    .A2(_01302_),
    .B1(_01896_),
    .B2(_02759_),
    .Y(_06091_)
  );
  sg13g2_a21oi_1 _16003_ (
    .A1(_07370_),
    .A2(_03954_),
    .B1(_00899_),
    .Y(_06092_)
  );
  sg13g2_nor4_1 _16004_ (
    .A(addr_i_8_),
    .B(_06090_),
    .C(_06091_),
    .D(_06092_),
    .Y(_06093_)
  );
  sg13g2_nand2_1 _16005_ (
    .A(_01527_),
    .B(_01588_),
    .Y(_06094_)
  );
  sg13g2_nand2_1 _16006_ (
    .A(addr_i_4_),
    .B(_00448_),
    .Y(_06095_)
  );
  sg13g2_a21oi_1 _16007_ (
    .A1(_01267_),
    .A2(_06095_),
    .B1(addr_i_3_),
    .Y(_06096_)
  );
  sg13g2_a22oi_1 _16008_ (
    .A1(addr_i_3_),
    .A2(_06094_),
    .B1(_06096_),
    .B2(_05452_),
    .Y(_06097_)
  );
  sg13g2_a21oi_1 _16009_ (
    .A1(_05856_),
    .A2(_06884_),
    .B1(_00014_),
    .Y(_06098_)
  );
  sg13g2_o21ai_1 _16010_ (
    .A1(addr_i_4_),
    .A2(_06098_),
    .B1(_00520_),
    .Y(_06100_)
  );
  sg13g2_o21ai_1 _16011_ (
    .A1(_02064_),
    .A2(_01339_),
    .B1(_01208_),
    .Y(_06101_)
  );
  sg13g2_nor2_1 _16012_ (
    .A(_05218_),
    .B(_00561_),
    .Y(_06102_)
  );
  sg13g2_a221oi_1 _16013_ (
    .A1(_01517_),
    .A2(_06100_),
    .B1(_06101_),
    .B2(addr_i_4_),
    .C1(_06102_),
    .Y(_06103_)
  );
  sg13g2_nor3_1 _16014_ (
    .A(_03242_),
    .B(_06097_),
    .C(_06103_),
    .Y(_06104_)
  );
  sg13g2_nor3_1 _16015_ (
    .A(_03073_),
    .B(_06093_),
    .C(_06104_),
    .Y(_06105_)
  );
  sg13g2_nor3_1 _16016_ (
    .A(addr_i_2_),
    .B(_01972_),
    .C(_03690_),
    .Y(_06106_)
  );
  sg13g2_a21oi_1 _16017_ (
    .A1(_00050_),
    .A2(_01441_),
    .B1(_00967_),
    .Y(_06107_)
  );
  sg13g2_a22oi_1 _16018_ (
    .A1(_02803_),
    .A2(_00686_),
    .B1(_06106_),
    .B2(_06107_),
    .Y(_06108_)
  );
  sg13g2_nand2_1 _16019_ (
    .A(_06895_),
    .B(_00943_),
    .Y(_06109_)
  );
  sg13g2_o21ai_1 _16020_ (
    .A1(_08100_),
    .A2(_03170_),
    .B1(addr_i_3_),
    .Y(_06111_)
  );
  sg13g2_a21oi_1 _16021_ (
    .A1(_00948_),
    .A2(_06111_),
    .B1(addr_i_4_),
    .Y(_06112_)
  );
  sg13g2_a22oi_1 _16022_ (
    .A1(addr_i_7_),
    .A2(_06109_),
    .B1(_06112_),
    .B2(_00629_),
    .Y(_06113_)
  );
  sg13g2_o21ai_1 _16023_ (
    .A1(addr_i_3_),
    .A2(_06108_),
    .B1(_06113_),
    .Y(_06114_)
  );
  sg13g2_nor2_1 _16024_ (
    .A(_08896_),
    .B(_07658_),
    .Y(_06115_)
  );
  sg13g2_o21ai_1 _16025_ (
    .A1(addr_i_3_),
    .A2(_06115_),
    .B1(_02001_),
    .Y(_06116_)
  );
  sg13g2_a21oi_1 _16026_ (
    .A1(_00520_),
    .A2(_06862_),
    .B1(_04461_),
    .Y(_06117_)
  );
  sg13g2_a21oi_1 _16027_ (
    .A1(_01527_),
    .A2(_03875_),
    .B1(addr_i_4_),
    .Y(_06118_)
  );
  sg13g2_a22oi_1 _16028_ (
    .A1(addr_i_4_),
    .A2(_06116_),
    .B1(_06117_),
    .B2(_06118_),
    .Y(_06119_)
  );
  sg13g2_nor2_1 _16029_ (
    .A(_00600_),
    .B(_06119_),
    .Y(_06120_)
  );
  sg13g2_o21ai_1 _16030_ (
    .A1(_02264_),
    .A2(_03106_),
    .B1(addr_i_3_),
    .Y(_06122_)
  );
  sg13g2_a21oi_1 _16031_ (
    .A1(_08708_),
    .A2(_02076_),
    .B1(_01420_),
    .Y(_06123_)
  );
  sg13g2_a21oi_1 _16032_ (
    .A1(_06122_),
    .A2(_06123_),
    .B1(_08830_),
    .Y(_06124_)
  );
  sg13g2_nor2_1 _16033_ (
    .A(_06120_),
    .B(_06124_),
    .Y(_06125_)
  );
  sg13g2_a21oi_1 _16034_ (
    .A1(_06114_),
    .A2(_06125_),
    .B1(_02221_),
    .Y(_06126_)
  );
  sg13g2_nand2_1 _16035_ (
    .A(_08796_),
    .B(_02052_),
    .Y(_06127_)
  );
  sg13g2_a22oi_1 _16036_ (
    .A1(addr_i_3_),
    .A2(_06127_),
    .B1(_00119_),
    .B2(addr_i_7_),
    .Y(_06128_)
  );
  sg13g2_nor2_1 _16037_ (
    .A(_07746_),
    .B(_01022_),
    .Y(_06129_)
  );
  sg13g2_nor2_1 _16038_ (
    .A(addr_i_3_),
    .B(_06129_),
    .Y(_06130_)
  );
  sg13g2_o21ai_1 _16039_ (
    .A1(_05300_),
    .A2(_06130_),
    .B1(addr_i_2_),
    .Y(_06131_)
  );
  sg13g2_o21ai_1 _16040_ (
    .A1(_02496_),
    .A2(_00226_),
    .B1(_01319_),
    .Y(_06133_)
  );
  sg13g2_nand2_1 _16041_ (
    .A(addr_i_8_),
    .B(_06133_),
    .Y(_06134_)
  );
  sg13g2_a21o_1 _16042_ (
    .A1(_06128_),
    .A2(_06131_),
    .B1(_06134_),
    .X(_06135_)
  );
  sg13g2_a21oi_1 _16043_ (
    .A1(addr_i_4_),
    .A2(_03021_),
    .B1(_00279_),
    .Y(_06136_)
  );
  sg13g2_nor2_1 _16044_ (
    .A(_00825_),
    .B(_06136_),
    .Y(_06137_)
  );
  sg13g2_a21oi_1 _16045_ (
    .A1(_01658_),
    .A2(_00284_),
    .B1(_00293_),
    .Y(_06138_)
  );
  sg13g2_a221oi_1 _16046_ (
    .A1(_09494_),
    .A2(_00808_),
    .B1(_01026_),
    .B2(addr_i_7_),
    .C1(_06138_),
    .Y(_06139_)
  );
  sg13g2_a22oi_1 _16047_ (
    .A1(_00065_),
    .A2(_00965_),
    .B1(_01514_),
    .B2(_00001_),
    .Y(_06140_)
  );
  sg13g2_nor3_1 _16048_ (
    .A(_08343_),
    .B(_00006_),
    .C(_01782_),
    .Y(_06141_)
  );
  sg13g2_a21oi_1 _16049_ (
    .A1(_00032_),
    .A2(_05083_),
    .B1(_00008_),
    .Y(_06142_)
  );
  sg13g2_nor4_1 _16050_ (
    .A(addr_i_8_),
    .B(_06140_),
    .C(_06141_),
    .D(_06142_),
    .Y(_06144_)
  );
  sg13g2_o21ai_1 _16051_ (
    .A1(_02530_),
    .A2(_06139_),
    .B1(_06144_),
    .Y(_06145_)
  );
  sg13g2_o21ai_1 _16052_ (
    .A1(_06135_),
    .A2(_06137_),
    .B1(_06145_),
    .Y(_06146_)
  );
  sg13g2_nand2_1 _16053_ (
    .A(_00545_),
    .B(_04421_),
    .Y(_06147_)
  );
  sg13g2_nor2_1 _16054_ (
    .A(_02471_),
    .B(_02076_),
    .Y(_06148_)
  );
  sg13g2_nor2_1 _16055_ (
    .A(_05856_),
    .B(_03139_),
    .Y(_06149_)
  );
  sg13g2_a22oi_1 _16056_ (
    .A1(_01888_),
    .A2(_02152_),
    .B1(_00304_),
    .B2(addr_i_3_),
    .Y(_06150_)
  );
  sg13g2_a22oi_1 _16057_ (
    .A1(_01768_),
    .A2(_06149_),
    .B1(_06150_),
    .B2(addr_i_7_),
    .Y(_06151_)
  );
  sg13g2_a22oi_1 _16058_ (
    .A1(_00578_),
    .A2(_06148_),
    .B1(_06151_),
    .B2(addr_i_8_),
    .Y(_06152_)
  );
  sg13g2_o21ai_1 _16059_ (
    .A1(_08896_),
    .A2(_00383_),
    .B1(addr_i_3_),
    .Y(_06153_)
  );
  sg13g2_nand3_1 _16060_ (
    .A(_01738_),
    .B(_03324_),
    .C(_06153_),
    .Y(_06155_)
  );
  sg13g2_o21ai_1 _16061_ (
    .A1(_00050_),
    .A2(_02470_),
    .B1(addr_i_8_),
    .Y(_06156_)
  );
  sg13g2_a221oi_1 _16062_ (
    .A1(addr_i_4_),
    .A2(_04214_),
    .B1(_06155_),
    .B2(addr_i_6_),
    .C1(_06156_),
    .Y(_06157_)
  );
  sg13g2_nor2_1 _16063_ (
    .A(_06152_),
    .B(_06157_),
    .Y(_06158_)
  );
  sg13g2_a22oi_1 _16064_ (
    .A1(_02501_),
    .A2(_06147_),
    .B1(_06158_),
    .B2(addr_i_9_),
    .Y(_06159_)
  );
  sg13g2_a22oi_1 _16065_ (
    .A1(addr_i_9_),
    .A2(_06146_),
    .B1(_06159_),
    .B2(addr_i_10_),
    .Y(_06160_)
  );
  sg13g2_nor4_1 _16066_ (
    .A(addr_i_11_),
    .B(_06105_),
    .C(_06126_),
    .D(_06160_),
    .Y(_06161_)
  );
  sg13g2_or3_1 _16067_ (
    .A(addr_i_12_),
    .B(_06085_),
    .C(_06161_),
    .X(_06162_)
  );
  sg13g2_o21ai_1 _16068_ (
    .A1(_05972_),
    .A2(_05996_),
    .B1(_06162_),
    .Y(data_o_26_)
  );
  sg13g2_o21ai_1 _16069_ (
    .A1(_01507_),
    .A2(_01194_),
    .B1(_01436_),
    .Y(_06163_)
  );
  sg13g2_nand3_1 _16070_ (
    .A(_00764_),
    .B(_03340_),
    .C(_06163_),
    .Y(_06166_)
  );
  sg13g2_a22oi_1 _16071_ (
    .A1(_01095_),
    .A2(_02592_),
    .B1(_06166_),
    .B2(addr_i_3_),
    .Y(_06167_)
  );
  sg13g2_nand3_1 _16072_ (
    .A(_01343_),
    .B(_01601_),
    .C(_01618_),
    .Y(_06168_)
  );
  sg13g2_a21oi_1 _16073_ (
    .A1(_01155_),
    .A2(_00930_),
    .B1(_01104_),
    .Y(_06169_)
  );
  sg13g2_a22oi_1 _16074_ (
    .A1(addr_i_4_),
    .A2(_06168_),
    .B1(_06169_),
    .B2(_00116_),
    .Y(_06170_)
  );
  sg13g2_o21ai_1 _16075_ (
    .A1(_06167_),
    .A2(_06170_),
    .B1(addr_i_8_),
    .Y(_06171_)
  );
  sg13g2_nand2_1 _16076_ (
    .A(_05599_),
    .B(_03445_),
    .Y(_06172_)
  );
  sg13g2_nor3_1 _16077_ (
    .A(_00098_),
    .B(_09498_),
    .C(_01020_),
    .Y(_06173_)
  );
  sg13g2_nor4_1 _16078_ (
    .A(addr_i_3_),
    .B(_01112_),
    .C(_02154_),
    .D(_01604_),
    .Y(_06174_)
  );
  sg13g2_a22oi_1 _16079_ (
    .A1(addr_i_3_),
    .A2(_06173_),
    .B1(_06174_),
    .B2(addr_i_4_),
    .Y(_06175_)
  );
  sg13g2_a22oi_1 _16080_ (
    .A1(_02257_),
    .A2(_06172_),
    .B1(_06175_),
    .B2(addr_i_8_),
    .Y(_06177_)
  );
  sg13g2_nor2_1 _16081_ (
    .A(addr_i_9_),
    .B(_06177_),
    .Y(_06178_)
  );
  sg13g2_a21oi_1 _16082_ (
    .A1(addr_i_4_),
    .A2(_08453_),
    .B1(addr_i_5_),
    .Y(_06179_)
  );
  sg13g2_o21ai_1 _16083_ (
    .A1(_01041_),
    .A2(_06179_),
    .B1(_01542_),
    .Y(_06180_)
  );
  sg13g2_o21ai_1 _16084_ (
    .A1(_02180_),
    .A2(_03450_),
    .B1(_00402_),
    .Y(_06181_)
  );
  sg13g2_o21ai_1 _16085_ (
    .A1(_01863_),
    .A2(_00746_),
    .B1(addr_i_4_),
    .Y(_06182_)
  );
  sg13g2_nand2b_1 _16086_ (
    .A_N(_04430_),
    .B(_06182_),
    .Y(_06183_)
  );
  sg13g2_a21oi_1 _16087_ (
    .A1(_05092_),
    .A2(_08022_),
    .B1(addr_i_2_),
    .Y(_06184_)
  );
  sg13g2_o21ai_1 _16088_ (
    .A1(_06183_),
    .A2(_06184_),
    .B1(addr_i_7_),
    .Y(_06185_)
  );
  sg13g2_nand4_1 _16089_ (
    .A(addr_i_8_),
    .B(_06180_),
    .C(_06181_),
    .D(_06185_),
    .Y(_06186_)
  );
  sg13g2_nand2_1 _16090_ (
    .A(_00545_),
    .B(_03871_),
    .Y(_06188_)
  );
  sg13g2_o21ai_1 _16091_ (
    .A1(_06220_),
    .A2(_01107_),
    .B1(addr_i_3_),
    .Y(_06189_)
  );
  sg13g2_a21oi_1 _16092_ (
    .A1(_02807_),
    .A2(_06189_),
    .B1(_02759_),
    .Y(_06190_)
  );
  sg13g2_a22oi_1 _16093_ (
    .A1(_01320_),
    .A2(_06188_),
    .B1(_06190_),
    .B2(addr_i_8_),
    .Y(_06191_)
  );
  sg13g2_a21oi_1 _16094_ (
    .A1(_00478_),
    .A2(_00940_),
    .B1(addr_i_4_),
    .Y(_06192_)
  );
  sg13g2_a22oi_1 _16095_ (
    .A1(_04022_),
    .A2(_00999_),
    .B1(_03565_),
    .B2(_06192_),
    .Y(_06193_)
  );
  sg13g2_or2_1 _16096_ (
    .A(addr_i_7_),
    .B(_06193_),
    .X(_06194_)
  );
  sg13g2_a21oi_1 _16097_ (
    .A1(_06191_),
    .A2(_06194_),
    .B1(_01351_),
    .Y(_06195_)
  );
  sg13g2_a221oi_1 _16098_ (
    .A1(_06171_),
    .A2(_06178_),
    .B1(_06186_),
    .B2(_06195_),
    .C1(_00511_),
    .Y(_06196_)
  );
  sg13g2_o21ai_1 _16099_ (
    .A1(_00347_),
    .A2(_01422_),
    .B1(_00731_),
    .Y(_06197_)
  );
  sg13g2_a21oi_1 _16100_ (
    .A1(_00872_),
    .A2(_03324_),
    .B1(_02777_),
    .Y(_06199_)
  );
  sg13g2_a22oi_1 _16101_ (
    .A1(addr_i_5_),
    .A2(_06197_),
    .B1(_06199_),
    .B2(_02171_),
    .Y(_06200_)
  );
  sg13g2_nor2_1 _16102_ (
    .A(_07403_),
    .B(_06200_),
    .Y(_06201_)
  );
  sg13g2_a21oi_1 _16103_ (
    .A1(addr_i_3_),
    .A2(_08553_),
    .B1(_00279_),
    .Y(_06202_)
  );
  sg13g2_nor2_1 _16104_ (
    .A(_00238_),
    .B(_01093_),
    .Y(_06203_)
  );
  sg13g2_a22oi_1 _16105_ (
    .A1(_02063_),
    .A2(_06203_),
    .B1(_00743_),
    .B2(addr_i_4_),
    .Y(_06204_)
  );
  sg13g2_a22oi_1 _16106_ (
    .A1(addr_i_4_),
    .A2(_06202_),
    .B1(_06204_),
    .B2(_00600_),
    .Y(_06205_)
  );
  sg13g2_nand2_1 _16107_ (
    .A(addr_i_2_),
    .B(_00713_),
    .Y(_06206_)
  );
  sg13g2_a22oi_1 _16108_ (
    .A1(_00822_),
    .A2(_01869_),
    .B1(_02731_),
    .B2(_01402_),
    .Y(_06207_)
  );
  sg13g2_o21ai_1 _16109_ (
    .A1(_01954_),
    .A2(_00746_),
    .B1(_01472_),
    .Y(_06208_)
  );
  sg13g2_o21ai_1 _16110_ (
    .A1(_08464_),
    .A2(_00514_),
    .B1(_06208_),
    .Y(_06210_)
  );
  sg13g2_a21oi_1 _16111_ (
    .A1(_00550_),
    .A2(_08941_),
    .B1(_00557_),
    .Y(_06211_)
  );
  sg13g2_nor4_1 _16112_ (
    .A(addr_i_2_),
    .B(_01011_),
    .C(_00319_),
    .D(_06211_),
    .Y(_06212_)
  );
  sg13g2_a21oi_1 _16113_ (
    .A1(_00276_),
    .A2(_06210_),
    .B1(_06212_),
    .Y(_06213_)
  );
  sg13g2_o21ai_1 _16114_ (
    .A1(_06206_),
    .A2(_06207_),
    .B1(_06213_),
    .Y(_06214_)
  );
  sg13g2_or3_1 _16115_ (
    .A(_06201_),
    .B(_06205_),
    .C(_06214_),
    .X(_06215_)
  );
  sg13g2_a21oi_1 _16116_ (
    .A1(_05070_),
    .A2(_00104_),
    .B1(_02387_),
    .Y(_06216_)
  );
  sg13g2_a21oi_1 _16117_ (
    .A1(_02404_),
    .A2(_01645_),
    .B1(_06216_),
    .Y(_06217_)
  );
  sg13g2_nand2_1 _16118_ (
    .A(_00017_),
    .B(_03854_),
    .Y(_06218_)
  );
  sg13g2_o21ai_1 _16119_ (
    .A1(addr_i_2_),
    .A2(_06217_),
    .B1(_06218_),
    .Y(_06219_)
  );
  sg13g2_o21ai_1 _16120_ (
    .A1(_00384_),
    .A2(_04483_),
    .B1(addr_i_3_),
    .Y(_06221_)
  );
  sg13g2_a21oi_1 _16121_ (
    .A1(_00646_),
    .A2(_06221_),
    .B1(addr_i_2_),
    .Y(_06222_)
  );
  sg13g2_nand2_1 _16122_ (
    .A(_08332_),
    .B(_00441_),
    .Y(_06223_)
  );
  sg13g2_a21oi_1 _16123_ (
    .A1(_03150_),
    .A2(_06223_),
    .B1(_02420_),
    .Y(_06224_)
  );
  sg13g2_a21oi_1 _16124_ (
    .A1(_00386_),
    .A2(_00644_),
    .B1(addr_i_8_),
    .Y(_06225_)
  );
  sg13g2_o21ai_1 _16125_ (
    .A1(addr_i_3_),
    .A2(_06224_),
    .B1(_06225_),
    .Y(_06226_)
  );
  sg13g2_a22oi_1 _16126_ (
    .A1(addr_i_6_),
    .A2(_06219_),
    .B1(_06222_),
    .B2(_06226_),
    .Y(_06227_)
  );
  sg13g2_nand2_1 _16127_ (
    .A(_00158_),
    .B(_07503_),
    .Y(_06228_)
  );
  sg13g2_o21ai_1 _16128_ (
    .A1(_00294_),
    .A2(_00010_),
    .B1(_00072_),
    .Y(_06229_)
  );
  sg13g2_nand3_1 _16129_ (
    .A(_06228_),
    .B(_02661_),
    .C(_06229_),
    .Y(_06230_)
  );
  sg13g2_nor2_1 _16130_ (
    .A(_00449_),
    .B(_02420_),
    .Y(_06232_)
  );
  sg13g2_nand2_1 _16131_ (
    .A(_00427_),
    .B(_06232_),
    .Y(_06233_)
  );
  sg13g2_nand2_1 _16132_ (
    .A(addr_i_8_),
    .B(_06784_),
    .Y(_06234_)
  );
  sg13g2_a221oi_1 _16133_ (
    .A1(_01324_),
    .A2(_06230_),
    .B1(_06233_),
    .B2(addr_i_3_),
    .C1(_06234_),
    .Y(_06235_)
  );
  sg13g2_nor3_1 _16134_ (
    .A(addr_i_9_),
    .B(_06227_),
    .C(_06235_),
    .Y(_06236_)
  );
  sg13g2_a22oi_1 _16135_ (
    .A1(addr_i_9_),
    .A2(_06215_),
    .B1(_06236_),
    .B2(addr_i_10_),
    .Y(_06237_)
  );
  sg13g2_nor3_1 _16136_ (
    .A(addr_i_11_),
    .B(_06196_),
    .C(_06237_),
    .Y(_06238_)
  );
  sg13g2_a21oi_1 _16137_ (
    .A1(_06228_),
    .A2(_06095_),
    .B1(addr_i_5_),
    .Y(_06239_)
  );
  sg13g2_a21oi_1 _16138_ (
    .A1(_01131_),
    .A2(_02626_),
    .B1(_00227_),
    .Y(_06240_)
  );
  sg13g2_o21ai_1 _16139_ (
    .A1(addr_i_3_),
    .A2(_06240_),
    .B1(_01533_),
    .Y(_06241_)
  );
  sg13g2_o21ai_1 _16140_ (
    .A1(_06239_),
    .A2(_06241_),
    .B1(_01119_),
    .Y(_06243_)
  );
  sg13g2_a21oi_1 _16141_ (
    .A1(_00938_),
    .A2(_01175_),
    .B1(addr_i_4_),
    .Y(_06244_)
  );
  sg13g2_a21oi_1 _16142_ (
    .A1(_01445_),
    .A2(_09226_),
    .B1(_06244_),
    .Y(_06245_)
  );
  sg13g2_o21ai_1 _16143_ (
    .A1(addr_i_3_),
    .A2(_06245_),
    .B1(_04808_),
    .Y(_06246_)
  );
  sg13g2_a22oi_1 _16144_ (
    .A1(_03927_),
    .A2(_02695_),
    .B1(addr_i_3_),
    .B2(_08830_),
    .Y(_06247_)
  );
  sg13g2_a22oi_1 _16145_ (
    .A1(_00440_),
    .A2(_06246_),
    .B1(_06247_),
    .B2(addr_i_9_),
    .Y(_06248_)
  );
  sg13g2_a22oi_1 _16146_ (
    .A1(_06243_),
    .A2(_06248_),
    .B1(addr_i_10_),
    .B2(_00781_),
    .Y(_06249_)
  );
  sg13g2_a21oi_1 _16147_ (
    .A1(_05645_),
    .A2(_00667_),
    .B1(_00808_),
    .Y(_06250_)
  );
  sg13g2_nor2_1 _16148_ (
    .A(_02040_),
    .B(_06250_),
    .Y(_06251_)
  );
  sg13g2_o21ai_1 _16149_ (
    .A1(_06249_),
    .A2(_06251_),
    .B1(addr_i_11_),
    .Y(_06252_)
  );
  sg13g2_nor2b_1 _16150_ (
    .A(_06238_),
    .B_N(_06252_),
    .Y(_06254_)
  );
  sg13g2_a21oi_1 _16151_ (
    .A1(_00764_),
    .A2(_01795_),
    .B1(_02796_),
    .Y(_06255_)
  );
  sg13g2_a22oi_1 _16152_ (
    .A1(_00223_),
    .A2(_02090_),
    .B1(_06255_),
    .B2(_01794_),
    .Y(_06256_)
  );
  sg13g2_nor2_1 _16153_ (
    .A(_00789_),
    .B(_02115_),
    .Y(_06257_)
  );
  sg13g2_a21oi_1 _16154_ (
    .A1(_03575_),
    .A2(_01199_),
    .B1(addr_i_3_),
    .Y(_06258_)
  );
  sg13g2_nor4_1 _16155_ (
    .A(addr_i_4_),
    .B(_08310_),
    .C(_06257_),
    .D(_06258_),
    .Y(_06259_)
  );
  sg13g2_o21ai_1 _16156_ (
    .A1(_06256_),
    .A2(_06259_),
    .B1(_01767_),
    .Y(_06260_)
  );
  sg13g2_a21oi_1 _16157_ (
    .A1(_00477_),
    .A2(_01175_),
    .B1(addr_i_3_),
    .Y(_06261_)
  );
  sg13g2_a21oi_1 _16158_ (
    .A1(_00155_),
    .A2(_04632_),
    .B1(addr_i_5_),
    .Y(_06262_)
  );
  sg13g2_o21ai_1 _16159_ (
    .A1(_06261_),
    .A2(_06262_),
    .B1(addr_i_4_),
    .Y(_06263_)
  );
  sg13g2_a21o_1 _16160_ (
    .A1(_00394_),
    .A2(_06263_),
    .B1(_01034_),
    .X(_06265_)
  );
  sg13g2_nand4_1 _16161_ (
    .A(addr_i_5_),
    .B(_02501_),
    .C(_00409_),
    .D(_01749_),
    .Y(_06266_)
  );
  sg13g2_a21oi_1 _16162_ (
    .A1(_00945_),
    .A2(_07503_),
    .B1(_01643_),
    .Y(_06267_)
  );
  sg13g2_nor2_1 _16163_ (
    .A(_01099_),
    .B(_06267_),
    .Y(_06268_)
  );
  sg13g2_a22oi_1 _16164_ (
    .A1(_00697_),
    .A2(_01872_),
    .B1(_03132_),
    .B2(addr_i_4_),
    .Y(_06269_)
  );
  sg13g2_a22oi_1 _16165_ (
    .A1(_00529_),
    .A2(_00850_),
    .B1(_06268_),
    .B2(_06269_),
    .Y(_06270_)
  );
  sg13g2_a21oi_1 _16166_ (
    .A1(_01125_),
    .A2(_00353_),
    .B1(addr_i_4_),
    .Y(_06271_)
  );
  sg13g2_o21ai_1 _16167_ (
    .A1(_02698_),
    .A2(_06271_),
    .B1(_00708_),
    .Y(_06272_)
  );
  sg13g2_nand4_1 _16168_ (
    .A(_06265_),
    .B(_06266_),
    .C(_06270_),
    .D(_06272_),
    .Y(_06273_)
  );
  sg13g2_o21ai_1 _16169_ (
    .A1(addr_i_7_),
    .A2(_05652_),
    .B1(_02956_),
    .Y(_06274_)
  );
  sg13g2_mux2_1 _16170_ (
    .A0(_01949_),
    .A1(_02405_),
    .S(addr_i_3_),
    .X(_06277_)
  );
  sg13g2_nor2_1 _16171_ (
    .A(addr_i_2_),
    .B(_00982_),
    .Y(_06278_)
  );
  sg13g2_a22oi_1 _16172_ (
    .A1(addr_i_2_),
    .A2(_06277_),
    .B1(_06278_),
    .B2(_01794_),
    .Y(_06279_)
  );
  sg13g2_a21oi_1 _16173_ (
    .A1(addr_i_3_),
    .A2(_06274_),
    .B1(_06279_),
    .Y(_06280_)
  );
  sg13g2_o21ai_1 _16174_ (
    .A1(_00807_),
    .A2(_06280_),
    .B1(_03029_),
    .Y(_06281_)
  );
  sg13g2_a221oi_1 _16175_ (
    .A1(_01613_),
    .A2(_06260_),
    .B1(_06273_),
    .B2(_05214_),
    .C1(_06281_),
    .Y(_06282_)
  );
  sg13g2_a22oi_1 _16176_ (
    .A1(_00617_),
    .A2(_04443_),
    .B1(_02374_),
    .B2(_00436_),
    .Y(_06283_)
  );
  sg13g2_nand2b_1 _16177_ (
    .A_N(_06283_),
    .B(addr_i_3_),
    .Y(_06284_)
  );
  sg13g2_nand2_1 _16178_ (
    .A(_05025_),
    .B(_02459_),
    .Y(_06285_)
  );
  sg13g2_o21ai_1 _16179_ (
    .A1(addr_i_3_),
    .A2(_01326_),
    .B1(_06285_),
    .Y(_06286_)
  );
  sg13g2_a21oi_1 _16180_ (
    .A1(_00016_),
    .A2(_01273_),
    .B1(addr_i_4_),
    .Y(_06288_)
  );
  sg13g2_o21ai_1 _16181_ (
    .A1(_03577_),
    .A2(_06288_),
    .B1(addr_i_3_),
    .Y(_06289_)
  );
  sg13g2_nand2b_1 _16182_ (
    .A_N(_06286_),
    .B(_06289_),
    .Y(_06290_)
  );
  sg13g2_a221oi_1 _16183_ (
    .A1(_00402_),
    .A2(_00031_),
    .B1(_06290_),
    .B2(addr_i_5_),
    .C1(addr_i_8_),
    .Y(_06291_)
  );
  sg13g2_o21ai_1 _16184_ (
    .A1(_02639_),
    .A2(_00132_),
    .B1(addr_i_5_),
    .Y(_06292_)
  );
  sg13g2_a21oi_1 _16185_ (
    .A1(_07879_),
    .A2(_07038_),
    .B1(addr_i_2_),
    .Y(_06293_)
  );
  sg13g2_a22oi_1 _16186_ (
    .A1(_01159_),
    .A2(_07879_),
    .B1(_02632_),
    .B2(_02287_),
    .Y(_06294_)
  );
  sg13g2_a22oi_1 _16187_ (
    .A1(_06292_),
    .A2(_06293_),
    .B1(_06294_),
    .B2(addr_i_3_),
    .Y(_06295_)
  );
  sg13g2_o21ai_1 _16188_ (
    .A1(_01587_),
    .A2(_01194_),
    .B1(addr_i_4_),
    .Y(_06296_)
  );
  sg13g2_o21ai_1 _16189_ (
    .A1(_00183_),
    .A2(_09495_),
    .B1(addr_i_2_),
    .Y(_06297_)
  );
  sg13g2_a21oi_1 _16190_ (
    .A1(_06296_),
    .A2(_06297_),
    .B1(_00531_),
    .Y(_06299_)
  );
  sg13g2_nor4_1 _16191_ (
    .A(_01043_),
    .B(_03587_),
    .C(_06295_),
    .D(_06299_),
    .Y(_06300_)
  );
  sg13g2_a22oi_1 _16192_ (
    .A1(_06284_),
    .A2(_06291_),
    .B1(_06300_),
    .B2(_09326_),
    .Y(_06301_)
  );
  sg13g2_a21oi_1 _16193_ (
    .A1(addr_i_2_),
    .A2(_01928_),
    .B1(_00497_),
    .Y(_06302_)
  );
  sg13g2_nor2_1 _16194_ (
    .A(addr_i_4_),
    .B(_06017_),
    .Y(_06303_)
  );
  sg13g2_o21ai_1 _16195_ (
    .A1(_01929_),
    .A2(_06303_),
    .B1(addr_i_3_),
    .Y(_06304_)
  );
  sg13g2_nand2_1 _16196_ (
    .A(_00342_),
    .B(_01920_),
    .Y(_06305_)
  );
  sg13g2_nand2_1 _16197_ (
    .A(addr_i_6_),
    .B(_01914_),
    .Y(_06306_)
  );
  sg13g2_a21o_1 _16198_ (
    .A1(_06305_),
    .A2(_06306_),
    .B1(addr_i_3_),
    .X(_06307_)
  );
  sg13g2_nand3_1 _16199_ (
    .A(_06302_),
    .B(_06304_),
    .C(_06307_),
    .Y(_06308_)
  );
  sg13g2_nand2_1 _16200_ (
    .A(addr_i_8_),
    .B(_04937_),
    .Y(_06310_)
  );
  sg13g2_a21oi_1 _16201_ (
    .A1(_06110_),
    .A2(_06310_),
    .B1(_03497_),
    .Y(_06311_)
  );
  sg13g2_nor2_1 _16202_ (
    .A(addr_i_7_),
    .B(_06311_),
    .Y(_06312_)
  );
  sg13g2_o21ai_1 _16203_ (
    .A1(_09494_),
    .A2(_01107_),
    .B1(addr_i_6_),
    .Y(_06313_)
  );
  sg13g2_a22oi_1 _16204_ (
    .A1(_00228_),
    .A2(_06313_),
    .B1(addr_i_3_),
    .B2(_01559_),
    .Y(_06314_)
  );
  sg13g2_o21ai_1 _16205_ (
    .A1(addr_i_5_),
    .A2(_02781_),
    .B1(_01933_),
    .Y(_06315_)
  );
  sg13g2_a22oi_1 _16206_ (
    .A1(_08155_),
    .A2(_06315_),
    .B1(_05102_),
    .B2(addr_i_3_),
    .Y(_06316_)
  );
  sg13g2_a221oi_1 _16207_ (
    .A1(addr_i_4_),
    .A2(_06408_),
    .B1(_01936_),
    .B2(addr_i_5_),
    .C1(_08752_),
    .Y(_06317_)
  );
  sg13g2_nor3_1 _16208_ (
    .A(_04191_),
    .B(_06316_),
    .C(_06317_),
    .Y(_06318_)
  );
  sg13g2_a22oi_1 _16209_ (
    .A1(_06331_),
    .A2(_00518_),
    .B1(_06314_),
    .B2(_06318_),
    .Y(_06319_)
  );
  sg13g2_a221oi_1 _16210_ (
    .A1(_06308_),
    .A2(_06312_),
    .B1(_06319_),
    .B2(addr_i_7_),
    .C1(addr_i_9_),
    .Y(_06321_)
  );
  sg13g2_o21ai_1 _16211_ (
    .A1(_06301_),
    .A2(_06321_),
    .B1(_01774_),
    .Y(_06322_)
  );
  sg13g2_nand2_1 _16212_ (
    .A(_06282_),
    .B(_06322_),
    .Y(_06323_)
  );
  sg13g2_nand2_1 _16213_ (
    .A(_00535_),
    .B(_07636_),
    .Y(_06324_)
  );
  sg13g2_nand2_1 _16214_ (
    .A(addr_i_3_),
    .B(_01026_),
    .Y(_06325_)
  );
  sg13g2_a21oi_1 _16215_ (
    .A1(_06324_),
    .A2(_06325_),
    .B1(addr_i_5_),
    .Y(_06326_)
  );
  sg13g2_or2_1 _16216_ (
    .A(_01286_),
    .B(_06326_),
    .X(_06327_)
  );
  sg13g2_a21oi_1 _16217_ (
    .A1(addr_i_3_),
    .A2(_03112_),
    .B1(_00278_),
    .Y(_06328_)
  );
  sg13g2_o21ai_1 _16218_ (
    .A1(_01653_),
    .A2(_05999_),
    .B1(addr_i_2_),
    .Y(_06329_)
  );
  sg13g2_o21ai_1 _16219_ (
    .A1(addr_i_4_),
    .A2(_06328_),
    .B1(_06329_),
    .Y(_06330_)
  );
  sg13g2_nor2_1 _16220_ (
    .A(_01015_),
    .B(_00416_),
    .Y(_06332_)
  );
  sg13g2_a22oi_1 _16221_ (
    .A1(_03281_),
    .A2(_02383_),
    .B1(_04225_),
    .B2(addr_i_3_),
    .Y(_06333_)
  );
  sg13g2_a21oi_1 _16222_ (
    .A1(addr_i_3_),
    .A2(_06332_),
    .B1(_06333_),
    .Y(_06334_)
  );
  sg13g2_a21oi_1 _16223_ (
    .A1(_00584_),
    .A2(_00671_),
    .B1(addr_i_5_),
    .Y(_06335_)
  );
  sg13g2_o21ai_1 _16224_ (
    .A1(_01049_),
    .A2(_06335_),
    .B1(addr_i_3_),
    .Y(_06336_)
  );
  sg13g2_o21ai_1 _16225_ (
    .A1(_01519_),
    .A2(_02165_),
    .B1(_06336_),
    .Y(_06337_)
  );
  sg13g2_mux4_1 _16226_ (
    .A0(_06327_),
    .A1(_06330_),
    .A2(_06334_),
    .A3(_06337_),
    .S0(_06905_),
    .S1(_00367_),
    .X(_06338_)
  );
  sg13g2_nand2_1 _16227_ (
    .A(addr_i_3_),
    .B(_00104_),
    .Y(_06339_)
  );
  sg13g2_nor2_1 _16228_ (
    .A(_06220_),
    .B(_01902_),
    .Y(_06340_)
  );
  sg13g2_a21oi_1 _16229_ (
    .A1(_06339_),
    .A2(_06340_),
    .B1(_06717_),
    .Y(_06341_)
  );
  sg13g2_nand2_1 _16230_ (
    .A(addr_i_2_),
    .B(_03391_),
    .Y(_06343_)
  );
  sg13g2_a22oi_1 _16231_ (
    .A1(addr_i_4_),
    .A2(_00665_),
    .B1(_00920_),
    .B2(addr_i_2_),
    .Y(_06344_)
  );
  sg13g2_nor2_1 _16232_ (
    .A(_00351_),
    .B(_06344_),
    .Y(_06345_)
  );
  sg13g2_o21ai_1 _16233_ (
    .A1(_06341_),
    .A2(_06343_),
    .B1(_06345_),
    .Y(_06346_)
  );
  sg13g2_nor2_1 _16234_ (
    .A(_05745_),
    .B(_00914_),
    .Y(_06347_)
  );
  sg13g2_o21ai_1 _16235_ (
    .A1(_06347_),
    .A2(_04578_),
    .B1(_09473_),
    .Y(_06348_)
  );
  sg13g2_o21ai_1 _16236_ (
    .A1(_00503_),
    .A2(_00829_),
    .B1(_09486_),
    .Y(_06349_)
  );
  sg13g2_and3_1 _16237_ (
    .A(addr_i_8_),
    .B(_06348_),
    .C(_06349_),
    .X(_06350_)
  );
  sg13g2_o21ai_1 _16238_ (
    .A1(addr_i_3_),
    .A2(_04579_),
    .B1(_03871_),
    .Y(_06351_)
  );
  sg13g2_a22oi_1 _16239_ (
    .A1(addr_i_3_),
    .A2(_04355_),
    .B1(_00551_),
    .B2(_00548_),
    .Y(_06352_)
  );
  sg13g2_a22oi_1 _16240_ (
    .A1(_09138_),
    .A2(_06351_),
    .B1(_06352_),
    .B2(addr_i_8_),
    .Y(_06354_)
  );
  sg13g2_a21oi_1 _16241_ (
    .A1(addr_i_3_),
    .A2(_05299_),
    .B1(_02143_),
    .Y(_06355_)
  );
  sg13g2_nor2_1 _16242_ (
    .A(addr_i_2_),
    .B(_06355_),
    .Y(_06356_)
  );
  sg13g2_o21ai_1 _16243_ (
    .A1(_04430_),
    .A2(_06356_),
    .B1(_00779_),
    .Y(_06357_)
  );
  sg13g2_a221oi_1 _16244_ (
    .A1(_06346_),
    .A2(_06350_),
    .B1(_06354_),
    .B2(_06357_),
    .C1(_00243_),
    .Y(_06358_)
  );
  sg13g2_a21oi_1 _16245_ (
    .A1(_00397_),
    .A2(_06338_),
    .B1(_06358_),
    .Y(_06359_)
  );
  sg13g2_nor2_1 _16246_ (
    .A(addr_i_5_),
    .B(_00098_),
    .Y(_06360_)
  );
  sg13g2_a21oi_1 _16247_ (
    .A1(_01543_),
    .A2(_04396_),
    .B1(_08388_),
    .Y(_06361_)
  );
  sg13g2_a21oi_1 _16248_ (
    .A1(_02294_),
    .A2(_00434_),
    .B1(addr_i_4_),
    .Y(_06362_)
  );
  sg13g2_nor4_1 _16249_ (
    .A(addr_i_3_),
    .B(_06360_),
    .C(_06361_),
    .D(_06362_),
    .Y(_06363_)
  );
  sg13g2_o21ai_1 _16250_ (
    .A1(_01585_),
    .A2(_00759_),
    .B1(addr_i_4_),
    .Y(_06365_)
  );
  sg13g2_nor2b_1 _16251_ (
    .A(_09479_),
    .B_N(_06365_),
    .Y(_06366_)
  );
  sg13g2_nor2b_1 _16252_ (
    .A(_03339_),
    .B_N(_02282_),
    .Y(_06367_)
  );
  sg13g2_o21ai_1 _16253_ (
    .A1(_06363_),
    .A2(_06366_),
    .B1(_06367_),
    .Y(_06368_)
  );
  sg13g2_o21ai_1 _16254_ (
    .A1(_02990_),
    .A2(_04371_),
    .B1(_03085_),
    .Y(_06369_)
  );
  sg13g2_nor3_1 _16255_ (
    .A(addr_i_5_),
    .B(_00408_),
    .C(_02395_),
    .Y(_06370_)
  );
  sg13g2_a22oi_1 _16256_ (
    .A1(addr_i_5_),
    .A2(_06369_),
    .B1(_06370_),
    .B2(addr_i_7_),
    .Y(_06371_)
  );
  sg13g2_nand3_1 _16257_ (
    .A(_00956_),
    .B(addr_i_2_),
    .C(_00915_),
    .Y(_06372_)
  );
  sg13g2_nand4_1 _16258_ (
    .A(addr_i_7_),
    .B(_01037_),
    .C(_06372_),
    .D(_03604_),
    .Y(_06373_)
  );
  sg13g2_nand3b_1 _16259_ (
    .A_N(_06371_),
    .B(_06373_),
    .C(addr_i_8_),
    .Y(_06374_)
  );
  sg13g2_nand3_1 _16260_ (
    .A(_09326_),
    .B(_06368_),
    .C(_06374_),
    .Y(_06376_)
  );
  sg13g2_o21ai_1 _16261_ (
    .A1(_02772_),
    .A2(_00282_),
    .B1(addr_i_4_),
    .Y(_06377_)
  );
  sg13g2_a21oi_1 _16262_ (
    .A1(addr_i_4_),
    .A2(_02470_),
    .B1(_00520_),
    .Y(_06378_)
  );
  sg13g2_nor4_1 _16263_ (
    .A(_07514_),
    .B(_00474_),
    .C(_02182_),
    .D(_06378_),
    .Y(_06379_)
  );
  sg13g2_nor2_1 _16264_ (
    .A(addr_i_3_),
    .B(_01049_),
    .Y(_06380_)
  );
  sg13g2_nor3_1 _16265_ (
    .A(_08752_),
    .B(_09359_),
    .C(_02042_),
    .Y(_06381_)
  );
  sg13g2_a22oi_1 _16266_ (
    .A1(_05012_),
    .A2(_06380_),
    .B1(_06381_),
    .B2(_08830_),
    .Y(_06382_)
  );
  sg13g2_a22oi_1 _16267_ (
    .A1(_06377_),
    .A2(_06379_),
    .B1(_06382_),
    .B2(_04705_),
    .Y(_06383_)
  );
  sg13g2_nand3_1 _16268_ (
    .A(addr_i_5_),
    .B(_00695_),
    .C(_03607_),
    .Y(_06384_)
  );
  sg13g2_o21ai_1 _16269_ (
    .A1(addr_i_3_),
    .A2(_00170_),
    .B1(addr_i_6_),
    .Y(_06385_)
  );
  sg13g2_nand3_1 _16270_ (
    .A(addr_i_3_),
    .B(_03465_),
    .C(_05898_),
    .Y(_06388_)
  );
  sg13g2_nand2b_1 _16271_ (
    .A_N(_06385_),
    .B(_06388_),
    .Y(_06389_)
  );
  sg13g2_a21oi_1 _16272_ (
    .A1(_06384_),
    .A2(_06389_),
    .B1(_03930_),
    .Y(_06390_)
  );
  sg13g2_a21oi_1 _16273_ (
    .A1(_09226_),
    .A2(_00170_),
    .B1(_00399_),
    .Y(_06391_)
  );
  sg13g2_nand3_1 _16274_ (
    .A(addr_i_8_),
    .B(_01445_),
    .C(_08553_),
    .Y(_06392_)
  );
  sg13g2_o21ai_1 _16275_ (
    .A1(addr_i_3_),
    .A2(_06391_),
    .B1(_06392_),
    .Y(_06393_)
  );
  sg13g2_o21ai_1 _16276_ (
    .A1(_06390_),
    .A2(_06393_),
    .B1(_06630_),
    .Y(_06394_)
  );
  sg13g2_a21oi_1 _16277_ (
    .A1(_06383_),
    .A2(_06394_),
    .B1(_01773_),
    .Y(_06395_)
  );
  sg13g2_a21oi_1 _16278_ (
    .A1(_06376_),
    .A2(_06395_),
    .B1(_03040_),
    .Y(_06396_)
  );
  sg13g2_o21ai_1 _16279_ (
    .A1(addr_i_10_),
    .A2(_06359_),
    .B1(_06396_),
    .Y(_06397_)
  );
  sg13g2_a21oi_1 _16280_ (
    .A1(_06323_),
    .A2(_06397_),
    .B1(addr_i_12_),
    .Y(_06399_)
  );
  sg13g2_a21oi_1 _16281_ (
    .A1(addr_i_12_),
    .A2(_06254_),
    .B1(_06399_),
    .Y(data_o_27_)
  );
  sg13g2_nor2_1 _16282_ (
    .A(_06017_),
    .B(_00852_),
    .Y(_06400_)
  );
  sg13g2_a21oi_1 _16283_ (
    .A1(_01937_),
    .A2(_06305_),
    .B1(addr_i_3_),
    .Y(_06401_)
  );
  sg13g2_o21ai_1 _16284_ (
    .A1(_06400_),
    .A2(_06401_),
    .B1(_08708_),
    .Y(_06402_)
  );
  sg13g2_nand3_1 _16285_ (
    .A(addr_i_3_),
    .B(_02020_),
    .C(_08520_),
    .Y(_06403_)
  );
  sg13g2_o21ai_1 _16286_ (
    .A1(_08796_),
    .A2(_01914_),
    .B1(_06403_),
    .Y(_06404_)
  );
  sg13g2_nor2_1 _16287_ (
    .A(addr_i_3_),
    .B(addr_i_8_),
    .Y(_06405_)
  );
  sg13g2_nand2_1 _16288_ (
    .A(_02152_),
    .B(_06405_),
    .Y(_06406_)
  );
  sg13g2_nand2_1 _16289_ (
    .A(_06320_),
    .B(_00210_),
    .Y(_06407_)
  );
  sg13g2_a21oi_1 _16290_ (
    .A1(_06406_),
    .A2(_06407_),
    .B1(_05302_),
    .Y(_06409_)
  );
  sg13g2_a21oi_1 _16291_ (
    .A1(addr_i_2_),
    .A2(_06404_),
    .B1(_06409_),
    .Y(_06410_)
  );
  sg13g2_a21oi_1 _16292_ (
    .A1(_06402_),
    .A2(_06410_),
    .B1(addr_i_7_),
    .Y(_06411_)
  );
  sg13g2_nand2_1 _16293_ (
    .A(addr_i_2_),
    .B(_01537_),
    .Y(_06412_)
  );
  sg13g2_nor2_1 _16294_ (
    .A(_00938_),
    .B(_06412_),
    .Y(_06413_)
  );
  sg13g2_nand2_1 _16295_ (
    .A(_01537_),
    .B(addr_i_5_),
    .Y(_06414_)
  );
  sg13g2_a21oi_1 _16296_ (
    .A1(_05139_),
    .A2(_06414_),
    .B1(addr_i_2_),
    .Y(_06415_)
  );
  sg13g2_o21ai_1 _16297_ (
    .A1(_06413_),
    .A2(_06415_),
    .B1(addr_i_4_),
    .Y(_06416_)
  );
  sg13g2_o21ai_1 _16298_ (
    .A1(_00120_),
    .A2(_06017_),
    .B1(_05977_),
    .Y(_06417_)
  );
  sg13g2_a221oi_1 _16299_ (
    .A1(_00145_),
    .A2(_01917_),
    .B1(_06417_),
    .B2(_00554_),
    .C1(_08752_),
    .Y(_06418_)
  );
  sg13g2_o21ai_1 _16300_ (
    .A1(_04063_),
    .A2(_06198_),
    .B1(_06412_),
    .Y(_06420_)
  );
  sg13g2_a221oi_1 _16301_ (
    .A1(_07647_),
    .A2(_05901_),
    .B1(_06420_),
    .B2(_00091_),
    .C1(addr_i_3_),
    .Y(_06421_)
  );
  sg13g2_a22oi_1 _16302_ (
    .A1(_06416_),
    .A2(_06418_),
    .B1(_06421_),
    .B2(_06905_),
    .Y(_06422_)
  );
  sg13g2_o21ai_1 _16303_ (
    .A1(_06411_),
    .A2(_06422_),
    .B1(addr_i_9_),
    .Y(_06423_)
  );
  sg13g2_a21oi_1 _16304_ (
    .A1(_01410_),
    .A2(_04475_),
    .B1(addr_i_3_),
    .Y(_06424_)
  );
  sg13g2_a22oi_1 _16305_ (
    .A1(_07647_),
    .A2(_01134_),
    .B1(_06424_),
    .B2(_03652_),
    .Y(_06425_)
  );
  sg13g2_a21o_1 _16306_ (
    .A1(_02343_),
    .A2(_02592_),
    .B1(_07171_),
    .X(_06426_)
  );
  sg13g2_a22oi_1 _16307_ (
    .A1(addr_i_3_),
    .A2(_06426_),
    .B1(_02361_),
    .B2(addr_i_4_),
    .Y(_06427_)
  );
  sg13g2_o21ai_1 _16308_ (
    .A1(_06425_),
    .A2(_06427_),
    .B1(addr_i_8_),
    .Y(_06428_)
  );
  sg13g2_a21oi_1 _16309_ (
    .A1(_01077_),
    .A2(_04632_),
    .B1(_04373_),
    .Y(_06429_)
  );
  sg13g2_o21ai_1 _16310_ (
    .A1(_04681_),
    .A2(_06429_),
    .B1(_00377_),
    .Y(_06431_)
  );
  sg13g2_a22oi_1 _16311_ (
    .A1(_03167_),
    .A2(_00498_),
    .B1(_02514_),
    .B2(_00103_),
    .Y(_06432_)
  );
  sg13g2_nor2_1 _16312_ (
    .A(addr_i_8_),
    .B(_06432_),
    .Y(_06433_)
  );
  sg13g2_a21oi_1 _16313_ (
    .A1(_06431_),
    .A2(_06433_),
    .B1(addr_i_9_),
    .Y(_06434_)
  );
  sg13g2_nand2_1 _16314_ (
    .A(_06428_),
    .B(_06434_),
    .Y(_06435_)
  );
  sg13g2_nand2_1 _16315_ (
    .A(_06423_),
    .B(_06435_),
    .Y(_06436_)
  );
  sg13g2_a21oi_1 _16316_ (
    .A1(addr_i_4_),
    .A2(_05361_),
    .B1(_04683_),
    .Y(_06437_)
  );
  sg13g2_o21ai_1 _16317_ (
    .A1(addr_i_7_),
    .A2(_06437_),
    .B1(_01414_),
    .Y(_06438_)
  );
  sg13g2_o21ai_1 _16318_ (
    .A1(_00624_),
    .A2(_05765_),
    .B1(addr_i_3_),
    .Y(_06439_)
  );
  sg13g2_a21oi_1 _16319_ (
    .A1(_03710_),
    .A2(_06439_),
    .B1(_01308_),
    .Y(_06440_)
  );
  sg13g2_a22oi_1 _16320_ (
    .A1(addr_i_6_),
    .A2(_06438_),
    .B1(_06440_),
    .B2(_05883_),
    .Y(_06442_)
  );
  sg13g2_a21oi_1 _16321_ (
    .A1(_01581_),
    .A2(_02089_),
    .B1(addr_i_2_),
    .Y(_06443_)
  );
  sg13g2_o21ai_1 _16322_ (
    .A1(_03643_),
    .A2(_06443_),
    .B1(_05302_),
    .Y(_06444_)
  );
  sg13g2_nor2_1 _16323_ (
    .A(addr_i_3_),
    .B(_04915_),
    .Y(_06445_)
  );
  sg13g2_nand2_1 _16324_ (
    .A(_02349_),
    .B(_04295_),
    .Y(_06446_)
  );
  sg13g2_a221oi_1 _16325_ (
    .A1(_07879_),
    .A2(_04443_),
    .B1(_06446_),
    .B2(addr_i_4_),
    .C1(_00046_),
    .Y(_06447_)
  );
  sg13g2_a21o_1 _16326_ (
    .A1(_06444_),
    .A2(_06445_),
    .B1(_06447_),
    .X(_06448_)
  );
  sg13g2_mux2_1 _16327_ (
    .A0(_06442_),
    .A1(_06448_),
    .S(addr_i_8_),
    .X(_06449_)
  );
  sg13g2_a21oi_1 _16328_ (
    .A1(_00785_),
    .A2(_01029_),
    .B1(_04981_),
    .Y(_06450_)
  );
  sg13g2_a22oi_1 _16329_ (
    .A1(_01571_),
    .A2(_03922_),
    .B1(_06450_),
    .B2(_03501_),
    .Y(_06451_)
  );
  sg13g2_nor2_1 _16330_ (
    .A(_00588_),
    .B(_06451_),
    .Y(_06453_)
  );
  sg13g2_nand2_1 _16331_ (
    .A(_02694_),
    .B(_00573_),
    .Y(_06454_)
  );
  sg13g2_a21oi_1 _16332_ (
    .A1(_02732_),
    .A2(_06372_),
    .B1(addr_i_3_),
    .Y(_06455_)
  );
  sg13g2_o21ai_1 _16333_ (
    .A1(_01896_),
    .A2(_09348_),
    .B1(addr_i_4_),
    .Y(_06456_)
  );
  sg13g2_nand3_1 _16334_ (
    .A(_01354_),
    .B(_00429_),
    .C(_06456_),
    .Y(_06457_)
  );
  sg13g2_a22oi_1 _16335_ (
    .A1(addr_i_3_),
    .A2(_06454_),
    .B1(_06455_),
    .B2(_06457_),
    .Y(_06458_)
  );
  sg13g2_o21ai_1 _16336_ (
    .A1(_00743_),
    .A2(_01015_),
    .B1(_01302_),
    .Y(_06459_)
  );
  sg13g2_o21ai_1 _16337_ (
    .A1(_01445_),
    .A2(_02500_),
    .B1(addr_i_6_),
    .Y(_06460_)
  );
  sg13g2_a21oi_1 _16338_ (
    .A1(_06459_),
    .A2(_06460_),
    .B1(_07403_),
    .Y(_06461_)
  );
  sg13g2_o21ai_1 _16339_ (
    .A1(addr_i_6_),
    .A2(_01888_),
    .B1(_00700_),
    .Y(_06462_)
  );
  sg13g2_nand3_1 _16340_ (
    .A(_00276_),
    .B(_01815_),
    .C(_06462_),
    .Y(_06464_)
  );
  sg13g2_o21ai_1 _16341_ (
    .A1(addr_i_5_),
    .A2(_03288_),
    .B1(addr_i_2_),
    .Y(_06465_)
  );
  sg13g2_a21oi_1 _16342_ (
    .A1(_01301_),
    .A2(_06465_),
    .B1(_03652_),
    .Y(_06466_)
  );
  sg13g2_o21ai_1 _16343_ (
    .A1(_06464_),
    .A2(_06466_),
    .B1(_01174_),
    .Y(_06467_)
  );
  sg13g2_nor4_1 _16344_ (
    .A(_06453_),
    .B(_06458_),
    .C(_06461_),
    .D(_06467_),
    .Y(_06468_)
  );
  sg13g2_a21oi_1 _16345_ (
    .A1(_05203_),
    .A2(_06449_),
    .B1(_06468_),
    .Y(_06469_)
  );
  sg13g2_o21ai_1 _16346_ (
    .A1(addr_i_10_),
    .A2(_06436_),
    .B1(_06469_),
    .Y(_06470_)
  );
  sg13g2_nand2_1 _16347_ (
    .A(_03270_),
    .B(_06408_),
    .Y(_06471_)
  );
  sg13g2_o21ai_1 _16348_ (
    .A1(_00120_),
    .A2(_06414_),
    .B1(_06471_),
    .Y(_06472_)
  );
  sg13g2_nand2_1 _16349_ (
    .A(addr_i_6_),
    .B(_04075_),
    .Y(_06473_)
  );
  sg13g2_a21oi_1 _16350_ (
    .A1(_01087_),
    .A2(_06473_),
    .B1(addr_i_8_),
    .Y(_06475_)
  );
  sg13g2_nor2_1 _16351_ (
    .A(_00938_),
    .B(_05902_),
    .Y(_06476_)
  );
  sg13g2_a22oi_1 _16352_ (
    .A1(addr_i_4_),
    .A2(_06472_),
    .B1(_06475_),
    .B2(_06476_),
    .Y(_06477_)
  );
  sg13g2_nor2_1 _16353_ (
    .A(_01920_),
    .B(_05112_),
    .Y(_06478_)
  );
  sg13g2_o21ai_1 _16354_ (
    .A1(addr_i_4_),
    .A2(_06478_),
    .B1(_01589_),
    .Y(_06479_)
  );
  sg13g2_a221oi_1 _16355_ (
    .A1(_00644_),
    .A2(_00170_),
    .B1(_06479_),
    .B2(addr_i_5_),
    .C1(_00822_),
    .Y(_06480_)
  );
  sg13g2_a21oi_1 _16356_ (
    .A1(_07149_),
    .A2(_06477_),
    .B1(_06480_),
    .Y(_06481_)
  );
  sg13g2_a22oi_1 _16357_ (
    .A1(_01365_),
    .A2(_06021_),
    .B1(_06481_),
    .B2(addr_i_7_),
    .Y(_06482_)
  );
  sg13g2_a22oi_1 _16358_ (
    .A1(_00783_),
    .A2(_05076_),
    .B1(_02010_),
    .B2(_02891_),
    .Y(_06483_)
  );
  sg13g2_a221oi_1 _16359_ (
    .A1(_04461_),
    .A2(_07359_),
    .B1(_05757_),
    .B2(addr_i_4_),
    .C1(addr_i_8_),
    .Y(_06484_)
  );
  sg13g2_a21oi_1 _16360_ (
    .A1(addr_i_8_),
    .A2(_06483_),
    .B1(_06484_),
    .Y(_06486_)
  );
  sg13g2_o21ai_1 _16361_ (
    .A1(_07647_),
    .A2(_01917_),
    .B1(_01131_),
    .Y(_06487_)
  );
  sg13g2_a22oi_1 _16362_ (
    .A1(_02287_),
    .A2(_01917_),
    .B1(_01024_),
    .B2(addr_i_3_),
    .Y(_06488_)
  );
  sg13g2_a22oi_1 _16363_ (
    .A1(addr_i_3_),
    .A2(_06487_),
    .B1(_06488_),
    .B2(addr_i_5_),
    .Y(_06489_)
  );
  sg13g2_nor3_1 _16364_ (
    .A(_00779_),
    .B(_06486_),
    .C(_06489_),
    .Y(_06490_)
  );
  sg13g2_o21ai_1 _16365_ (
    .A1(_06482_),
    .A2(_06490_),
    .B1(addr_i_9_),
    .Y(_06491_)
  );
  sg13g2_a21oi_1 _16366_ (
    .A1(addr_i_2_),
    .A2(_04042_),
    .B1(_02265_),
    .Y(_06492_)
  );
  sg13g2_nor2_1 _16367_ (
    .A(_02530_),
    .B(_06492_),
    .Y(_06493_)
  );
  sg13g2_o21ai_1 _16368_ (
    .A1(_04679_),
    .A2(_06493_),
    .B1(_01861_),
    .Y(_06494_)
  );
  sg13g2_o21ai_1 _16369_ (
    .A1(_00252_),
    .A2(_00175_),
    .B1(addr_i_3_),
    .Y(_06495_)
  );
  sg13g2_a21oi_1 _16370_ (
    .A1(_09475_),
    .A2(_06495_),
    .B1(addr_i_6_),
    .Y(_06498_)
  );
  sg13g2_o21ai_1 _16371_ (
    .A1(_06519_),
    .A2(_06498_),
    .B1(_00276_),
    .Y(_06499_)
  );
  sg13g2_a22oi_1 _16372_ (
    .A1(addr_i_4_),
    .A2(_03545_),
    .B1(_01106_),
    .B2(_01276_),
    .Y(_06500_)
  );
  sg13g2_nor2_1 _16373_ (
    .A(_01757_),
    .B(_00521_),
    .Y(_06501_)
  );
  sg13g2_o21ai_1 _16374_ (
    .A1(_00011_),
    .A2(_06501_),
    .B1(addr_i_2_),
    .Y(_06502_)
  );
  sg13g2_o21ai_1 _16375_ (
    .A1(_00046_),
    .A2(_06500_),
    .B1(_06502_),
    .Y(_06503_)
  );
  sg13g2_a22oi_1 _16376_ (
    .A1(addr_i_6_),
    .A2(_00464_),
    .B1(_01659_),
    .B2(_00479_),
    .Y(_06504_)
  );
  sg13g2_a22oi_1 _16377_ (
    .A1(_00846_),
    .A2(_02942_),
    .B1(_06504_),
    .B2(_01494_),
    .Y(_06505_)
  );
  sg13g2_a21oi_1 _16378_ (
    .A1(_00429_),
    .A2(_06503_),
    .B1(_06505_),
    .Y(_06506_)
  );
  sg13g2_and3_1 _16379_ (
    .A(_09315_),
    .B(_06499_),
    .C(_06506_),
    .X(_06507_)
  );
  sg13g2_a21oi_1 _16380_ (
    .A1(_06494_),
    .A2(_06507_),
    .B1(addr_i_10_),
    .Y(_06509_)
  );
  sg13g2_nor2_1 _16381_ (
    .A(addr_i_3_),
    .B(_05925_),
    .Y(_06510_)
  );
  sg13g2_a21oi_1 _16382_ (
    .A1(addr_i_3_),
    .A2(_02517_),
    .B1(_00257_),
    .Y(_06511_)
  );
  sg13g2_o21ai_1 _16383_ (
    .A1(addr_i_4_),
    .A2(_06511_),
    .B1(_03346_),
    .Y(_06512_)
  );
  sg13g2_o21ai_1 _16384_ (
    .A1(_06510_),
    .A2(_06512_),
    .B1(_01324_),
    .Y(_06513_)
  );
  sg13g2_nor2_1 _16385_ (
    .A(_01014_),
    .B(_00789_),
    .Y(_06514_)
  );
  sg13g2_a21oi_1 _16386_ (
    .A1(_04981_),
    .A2(_01486_),
    .B1(_06514_),
    .Y(_06515_)
  );
  sg13g2_o21ai_1 _16387_ (
    .A1(_07215_),
    .A2(_01560_),
    .B1(_02404_),
    .Y(_06516_)
  );
  sg13g2_o21ai_1 _16388_ (
    .A1(_03652_),
    .A2(_06515_),
    .B1(_06516_),
    .Y(_06517_)
  );
  sg13g2_nor3_1 _16389_ (
    .A(_00342_),
    .B(_00586_),
    .C(_00025_),
    .Y(_06518_)
  );
  sg13g2_a22oi_1 _16390_ (
    .A1(addr_i_5_),
    .A2(_06517_),
    .B1(_06518_),
    .B2(addr_i_8_),
    .Y(_06520_)
  );
  sg13g2_a21oi_1 _16391_ (
    .A1(_03820_),
    .A2(_02898_),
    .B1(addr_i_3_),
    .Y(_06521_)
  );
  sg13g2_o21ai_1 _16392_ (
    .A1(_02203_),
    .A2(_06521_),
    .B1(_08011_),
    .Y(_06522_)
  );
  sg13g2_a21oi_1 _16393_ (
    .A1(_00381_),
    .A2(_01438_),
    .B1(_00190_),
    .Y(_06523_)
  );
  sg13g2_a21oi_1 _16394_ (
    .A1(_03497_),
    .A2(_02987_),
    .B1(_02344_),
    .Y(_06524_)
  );
  sg13g2_nor2_1 _16395_ (
    .A(_06523_),
    .B(_06524_),
    .Y(_06525_)
  );
  sg13g2_nand3_1 _16396_ (
    .A(_02405_),
    .B(_06522_),
    .C(_06525_),
    .Y(_06526_)
  );
  sg13g2_nand2_1 _16397_ (
    .A(addr_i_5_),
    .B(_00358_),
    .Y(_06527_)
  );
  sg13g2_nand2_1 _16398_ (
    .A(addr_i_3_),
    .B(_03545_),
    .Y(_06528_)
  );
  sg13g2_o21ai_1 _16399_ (
    .A1(_03919_),
    .A2(_03288_),
    .B1(_04373_),
    .Y(_06529_)
  );
  sg13g2_nand2_1 _16400_ (
    .A(_06528_),
    .B(_06529_),
    .Y(_06531_)
  );
  sg13g2_a22oi_1 _16401_ (
    .A1(addr_i_4_),
    .A2(_06527_),
    .B1(_06531_),
    .B2(_02405_),
    .Y(_06532_)
  );
  sg13g2_nor2_1 _16402_ (
    .A(_00782_),
    .B(_06532_),
    .Y(_06533_)
  );
  sg13g2_a221oi_1 _16403_ (
    .A1(_06513_),
    .A2(_06520_),
    .B1(_06526_),
    .B2(_06533_),
    .C1(_00925_),
    .Y(_06534_)
  );
  sg13g2_a21oi_1 _16404_ (
    .A1(_03540_),
    .A2(_05036_),
    .B1(addr_i_3_),
    .Y(_06535_)
  );
  sg13g2_nand2_1 _16405_ (
    .A(_00186_),
    .B(_00763_),
    .Y(_06536_)
  );
  sg13g2_o21ai_1 _16406_ (
    .A1(_06535_),
    .A2(_06536_),
    .B1(addr_i_4_),
    .Y(_06537_)
  );
  sg13g2_o21ai_1 _16407_ (
    .A1(addr_i_3_),
    .A2(_02638_),
    .B1(_01203_),
    .Y(_06538_)
  );
  sg13g2_nand2_1 _16408_ (
    .A(_00122_),
    .B(_06538_),
    .Y(_06539_)
  );
  sg13g2_nand3b_1 _16409_ (
    .A_N(_02622_),
    .B(_06537_),
    .C(_06539_),
    .Y(_06540_)
  );
  sg13g2_nand3_1 _16410_ (
    .A(_00262_),
    .B(_02297_),
    .C(_00719_),
    .Y(_06542_)
  );
  sg13g2_o21ai_1 _16411_ (
    .A1(_01850_),
    .A2(_06542_),
    .B1(_00629_),
    .Y(_06543_)
  );
  sg13g2_o21ai_1 _16412_ (
    .A1(_01445_),
    .A2(_09094_),
    .B1(addr_i_3_),
    .Y(_06544_)
  );
  sg13g2_a21oi_1 _16413_ (
    .A1(_04222_),
    .A2(_06544_),
    .B1(_00230_),
    .Y(_06545_)
  );
  sg13g2_a22oi_1 _16414_ (
    .A1(addr_i_6_),
    .A2(_06540_),
    .B1(_06543_),
    .B2(_06545_),
    .Y(_06546_)
  );
  sg13g2_a21oi_1 _16415_ (
    .A1(_00716_),
    .A2(_03660_),
    .B1(_08000_),
    .Y(_06547_)
  );
  sg13g2_o21ai_1 _16416_ (
    .A1(_00607_),
    .A2(_06547_),
    .B1(_01878_),
    .Y(_06548_)
  );
  sg13g2_a21o_1 _16417_ (
    .A1(_07072_),
    .A2(_02810_),
    .B1(_01103_),
    .X(_06549_)
  );
  sg13g2_o21ai_1 _16418_ (
    .A1(_00252_),
    .A2(_00303_),
    .B1(_01244_),
    .Y(_06550_)
  );
  sg13g2_nand3_1 _16419_ (
    .A(_04451_),
    .B(_02187_),
    .C(_06550_),
    .Y(_06551_)
  );
  sg13g2_nand2_1 _16420_ (
    .A(_04151_),
    .B(_07636_),
    .Y(_06553_)
  );
  sg13g2_o21ai_1 _16421_ (
    .A1(_00383_),
    .A2(_04849_),
    .B1(addr_i_3_),
    .Y(_06554_)
  );
  sg13g2_a21oi_1 _16422_ (
    .A1(_06553_),
    .A2(_06554_),
    .B1(addr_i_5_),
    .Y(_06555_)
  );
  sg13g2_a21oi_1 _16423_ (
    .A1(addr_i_7_),
    .A2(_06551_),
    .B1(_06555_),
    .Y(_06556_)
  );
  sg13g2_nand4_1 _16424_ (
    .A(addr_i_8_),
    .B(_06548_),
    .C(_06549_),
    .D(_06556_),
    .Y(_06557_)
  );
  sg13g2_nand2_1 _16425_ (
    .A(_01174_),
    .B(_06557_),
    .Y(_06558_)
  );
  sg13g2_o21ai_1 _16426_ (
    .A1(_06546_),
    .A2(_06558_),
    .B1(addr_i_11_),
    .Y(_06559_)
  );
  sg13g2_a22oi_1 _16427_ (
    .A1(_06491_),
    .A2(_06509_),
    .B1(_06534_),
    .B2(_06559_),
    .Y(_06560_)
  );
  sg13g2_a22oi_1 _16428_ (
    .A1(_03051_),
    .A2(_06470_),
    .B1(_06560_),
    .B2(addr_i_12_),
    .Y(_06561_)
  );
  sg13g2_a21o_1 _16429_ (
    .A1(_01892_),
    .A2(_04130_),
    .B1(_01357_),
    .X(_06562_)
  );
  sg13g2_o21ai_1 _16430_ (
    .A1(_06276_),
    .A2(_01732_),
    .B1(addr_i_4_),
    .Y(_06564_)
  );
  sg13g2_a21oi_1 _16431_ (
    .A1(_00677_),
    .A2(_06564_),
    .B1(_01935_),
    .Y(_06565_)
  );
  sg13g2_a21oi_1 _16432_ (
    .A1(_00516_),
    .A2(_01222_),
    .B1(addr_i_2_),
    .Y(_06566_)
  );
  sg13g2_a21oi_1 _16433_ (
    .A1(_00322_),
    .A2(_00074_),
    .B1(_06566_),
    .Y(_06567_)
  );
  sg13g2_o21ai_1 _16434_ (
    .A1(addr_i_7_),
    .A2(_02171_),
    .B1(_00949_),
    .Y(_06568_)
  );
  sg13g2_o21ai_1 _16435_ (
    .A1(addr_i_4_),
    .A2(_06567_),
    .B1(_06568_),
    .Y(_06569_)
  );
  sg13g2_o21ai_1 _16436_ (
    .A1(_06565_),
    .A2(_06569_),
    .B1(addr_i_8_),
    .Y(_06570_)
  );
  sg13g2_o21ai_1 _16437_ (
    .A1(addr_i_2_),
    .A2(_03139_),
    .B1(addr_i_3_),
    .Y(_06571_)
  );
  sg13g2_a21o_1 _16438_ (
    .A1(_00477_),
    .A2(_06571_),
    .B1(addr_i_5_),
    .X(_06572_)
  );
  sg13g2_o21ai_1 _16439_ (
    .A1(addr_i_3_),
    .A2(_05558_),
    .B1(_06572_),
    .Y(_06573_)
  );
  sg13g2_nor3_1 _16440_ (
    .A(addr_i_2_),
    .B(_00151_),
    .C(_01571_),
    .Y(_06575_)
  );
  sg13g2_a22oi_1 _16441_ (
    .A1(addr_i_2_),
    .A2(_00151_),
    .B1(_00600_),
    .B2(_06575_),
    .Y(_06576_)
  );
  sg13g2_a22oi_1 _16442_ (
    .A1(_00610_),
    .A2(_06573_),
    .B1(_06576_),
    .B2(addr_i_9_),
    .Y(_06577_)
  );
  sg13g2_a21oi_1 _16443_ (
    .A1(_00791_),
    .A2(_01285_),
    .B1(addr_i_5_),
    .Y(_06578_)
  );
  sg13g2_a22oi_1 _16444_ (
    .A1(addr_i_5_),
    .A2(_01633_),
    .B1(_01360_),
    .B2(_06578_),
    .Y(_06579_)
  );
  sg13g2_o21ai_1 _16445_ (
    .A1(_04705_),
    .A2(_06579_),
    .B1(_03731_),
    .Y(_06580_)
  );
  sg13g2_a21oi_1 _16446_ (
    .A1(_06570_),
    .A2(_06577_),
    .B1(_06580_),
    .Y(_06581_)
  );
  sg13g2_a22oi_1 _16447_ (
    .A1(_01350_),
    .A2(_06562_),
    .B1(_06581_),
    .B2(_01640_),
    .Y(_06582_)
  );
  sg13g2_a22oi_1 _16448_ (
    .A1(addr_i_2_),
    .A2(_05927_),
    .B1(_08188_),
    .B2(addr_i_5_),
    .Y(_06583_)
  );
  sg13g2_a22oi_1 _16449_ (
    .A1(_07116_),
    .A2(_01294_),
    .B1(_06583_),
    .B2(addr_i_3_),
    .Y(_06584_)
  );
  sg13g2_nor3_1 _16450_ (
    .A(_00294_),
    .B(_08941_),
    .C(_03110_),
    .Y(_06586_)
  );
  sg13g2_a22oi_1 _16451_ (
    .A1(_05634_),
    .A2(_01464_),
    .B1(_06586_),
    .B2(_06684_),
    .Y(_06587_)
  );
  sg13g2_o21ai_1 _16452_ (
    .A1(_09506_),
    .A2(_04176_),
    .B1(_08388_),
    .Y(_06588_)
  );
  sg13g2_nand2_1 _16453_ (
    .A(_06587_),
    .B(_06588_),
    .Y(_06589_)
  );
  sg13g2_o21ai_1 _16454_ (
    .A1(addr_i_3_),
    .A2(_03766_),
    .B1(_01406_),
    .Y(_06590_)
  );
  sg13g2_nor3_1 _16455_ (
    .A(_06298_),
    .B(_05910_),
    .C(_01244_),
    .Y(_06591_)
  );
  sg13g2_a21oi_1 _16456_ (
    .A1(addr_i_4_),
    .A2(_06590_),
    .B1(_06591_),
    .Y(_06592_)
  );
  sg13g2_o21ai_1 _16457_ (
    .A1(_03765_),
    .A2(_03194_),
    .B1(_05700_),
    .Y(_06593_)
  );
  sg13g2_nand3_1 _16458_ (
    .A(_04318_),
    .B(_01398_),
    .C(_06593_),
    .Y(_06594_)
  );
  sg13g2_nand2b_1 _16459_ (
    .A_N(_00493_),
    .B(_04933_),
    .Y(_06595_)
  );
  sg13g2_a221oi_1 _16460_ (
    .A1(_01319_),
    .A2(_06594_),
    .B1(_06595_),
    .B2(_09127_),
    .C1(addr_i_8_),
    .Y(_06597_)
  );
  sg13g2_o21ai_1 _16461_ (
    .A1(addr_i_7_),
    .A2(_06592_),
    .B1(_06597_),
    .Y(_06598_)
  );
  sg13g2_o21ai_1 _16462_ (
    .A1(_06584_),
    .A2(_06589_),
    .B1(_06598_),
    .Y(_06599_)
  );
  sg13g2_nor2_1 _16463_ (
    .A(_00715_),
    .B(_01097_),
    .Y(_06600_)
  );
  sg13g2_o21ai_1 _16464_ (
    .A1(_03132_),
    .A2(_04145_),
    .B1(_00385_),
    .Y(_06601_)
  );
  sg13g2_a21oi_1 _16465_ (
    .A1(_02578_),
    .A2(_06600_),
    .B1(_06601_),
    .Y(_06602_)
  );
  sg13g2_nand2_1 _16466_ (
    .A(_01837_),
    .B(_00960_),
    .Y(_06603_)
  );
  sg13g2_o21ai_1 _16467_ (
    .A1(addr_i_2_),
    .A2(_05297_),
    .B1(_06603_),
    .Y(_06604_)
  );
  sg13g2_nor2_1 _16468_ (
    .A(_00030_),
    .B(_00448_),
    .Y(_06605_)
  );
  sg13g2_o21ai_1 _16469_ (
    .A1(_01825_),
    .A2(_06605_),
    .B1(addr_i_5_),
    .Y(_06606_)
  );
  sg13g2_a21oi_1 _16470_ (
    .A1(_00211_),
    .A2(_00358_),
    .B1(addr_i_4_),
    .Y(_06609_)
  );
  sg13g2_a22oi_1 _16471_ (
    .A1(_06054_),
    .A2(_01044_),
    .B1(_06609_),
    .B2(addr_i_7_),
    .Y(_06610_)
  );
  sg13g2_a22oi_1 _16472_ (
    .A1(addr_i_7_),
    .A2(_06606_),
    .B1(_06610_),
    .B2(addr_i_8_),
    .Y(_06611_)
  );
  sg13g2_a21oi_1 _16473_ (
    .A1(_01118_),
    .A2(_06604_),
    .B1(_06611_),
    .Y(_06612_)
  );
  sg13g2_a221oi_1 _16474_ (
    .A1(addr_i_9_),
    .A2(_06599_),
    .B1(_06602_),
    .B2(_06612_),
    .C1(addr_i_10_),
    .Y(_06613_)
  );
  sg13g2_nand2_1 _16475_ (
    .A(_03853_),
    .B(_00712_),
    .Y(_06614_)
  );
  sg13g2_a21o_1 _16476_ (
    .A1(_05720_),
    .A2(_06614_),
    .B1(_00899_),
    .X(_06615_)
  );
  sg13g2_o21ai_1 _16477_ (
    .A1(_01160_),
    .A2(_00607_),
    .B1(_01460_),
    .Y(_06616_)
  );
  sg13g2_o21ai_1 _16478_ (
    .A1(_02427_),
    .A2(_02928_),
    .B1(addr_i_8_),
    .Y(_06617_)
  );
  sg13g2_nand2_1 _16479_ (
    .A(_00582_),
    .B(_00408_),
    .Y(_06618_)
  );
  sg13g2_a21oi_1 _16480_ (
    .A1(_01125_),
    .A2(_00762_),
    .B1(_01528_),
    .Y(_06620_)
  );
  sg13g2_a22oi_1 _16481_ (
    .A1(_00060_),
    .A2(_06618_),
    .B1(_06620_),
    .B2(_00324_),
    .Y(_06621_)
  );
  sg13g2_a22oi_1 _16482_ (
    .A1(_01542_),
    .A2(_06616_),
    .B1(_06617_),
    .B2(_06621_),
    .Y(_06622_)
  );
  sg13g2_a21oi_1 _16483_ (
    .A1(_00443_),
    .A2(_03445_),
    .B1(_00317_),
    .Y(_06623_)
  );
  sg13g2_a22oi_1 _16484_ (
    .A1(_00023_),
    .A2(_01309_),
    .B1(_06623_),
    .B2(addr_i_8_),
    .Y(_06624_)
  );
  sg13g2_nand2_1 _16485_ (
    .A(_06132_),
    .B(_00861_),
    .Y(_06625_)
  );
  sg13g2_a21oi_1 _16486_ (
    .A1(_06228_),
    .A2(_06625_),
    .B1(_00497_),
    .Y(_06626_)
  );
  sg13g2_o21ai_1 _16487_ (
    .A1(_06347_),
    .A2(_06626_),
    .B1(addr_i_7_),
    .Y(_06627_)
  );
  sg13g2_a221oi_1 _16488_ (
    .A1(_06615_),
    .A2(_06622_),
    .B1(_06624_),
    .B2(_06627_),
    .C1(_06652_),
    .Y(_06628_)
  );
  sg13g2_nand3_1 _16489_ (
    .A(_00554_),
    .B(_01672_),
    .C(_01199_),
    .Y(_06629_)
  );
  sg13g2_nand3_1 _16490_ (
    .A(addr_i_4_),
    .B(_01738_),
    .C(_00618_),
    .Y(_06631_)
  );
  sg13g2_a21oi_1 _16491_ (
    .A1(_06629_),
    .A2(_06631_),
    .B1(addr_i_5_),
    .Y(_06632_)
  );
  sg13g2_a22oi_1 _16492_ (
    .A1(_00967_),
    .A2(_05046_),
    .B1(_08410_),
    .B2(_03263_),
    .Y(_06633_)
  );
  sg13g2_o21ai_1 _16493_ (
    .A1(_06632_),
    .A2(_06633_),
    .B1(addr_i_3_),
    .Y(_06634_)
  );
  sg13g2_o21ai_1 _16494_ (
    .A1(_03919_),
    .A2(_00574_),
    .B1(_00228_),
    .Y(_06635_)
  );
  sg13g2_a22oi_1 _16495_ (
    .A1(addr_i_7_),
    .A2(_06635_),
    .B1(_01231_),
    .B2(addr_i_3_),
    .Y(_06636_)
  );
  sg13g2_nor2_1 _16496_ (
    .A(addr_i_8_),
    .B(_06636_),
    .Y(_06637_)
  );
  sg13g2_a22oi_1 _16497_ (
    .A1(_03809_),
    .A2(_00915_),
    .B1(_05280_),
    .B2(addr_i_2_),
    .Y(_06638_)
  );
  sg13g2_a21oi_1 _16498_ (
    .A1(_00050_),
    .A2(_02626_),
    .B1(_06638_),
    .Y(_06639_)
  );
  sg13g2_a21oi_1 _16499_ (
    .A1(_01527_),
    .A2(_00870_),
    .B1(_00007_),
    .Y(_06640_)
  );
  sg13g2_a21oi_1 _16500_ (
    .A1(addr_i_3_),
    .A2(_06639_),
    .B1(_06640_),
    .Y(_06642_)
  );
  sg13g2_nand2_1 _16501_ (
    .A(_09371_),
    .B(_02283_),
    .Y(_06643_)
  );
  sg13g2_a21o_1 _16502_ (
    .A1(_01067_),
    .A2(_06643_),
    .B1(_00100_),
    .X(_06644_)
  );
  sg13g2_nor2_1 _16503_ (
    .A(_02012_),
    .B(_02833_),
    .Y(_06645_)
  );
  sg13g2_o21ai_1 _16504_ (
    .A1(_02076_),
    .A2(_01222_),
    .B1(_01114_),
    .Y(_06646_)
  );
  sg13g2_a22oi_1 _16505_ (
    .A1(_03263_),
    .A2(_06644_),
    .B1(_06645_),
    .B2(_06646_),
    .Y(_06647_)
  );
  sg13g2_a22oi_1 _16506_ (
    .A1(addr_i_4_),
    .A2(_06642_),
    .B1(_06647_),
    .B2(_00782_),
    .Y(_06648_)
  );
  sg13g2_a21oi_1 _16507_ (
    .A1(_06634_),
    .A2(_06637_),
    .B1(_06648_),
    .Y(_06649_)
  );
  sg13g2_nor2_1 _16508_ (
    .A(_02221_),
    .B(_06649_),
    .Y(_06650_)
  );
  sg13g2_nor4_1 _16509_ (
    .A(addr_i_11_),
    .B(_06613_),
    .C(_06628_),
    .D(_06650_),
    .Y(_06651_)
  );
  sg13g2_nor3_1 _16510_ (
    .A(_00812_),
    .B(_06582_),
    .C(_06651_),
    .Y(_06653_)
  );
  sg13g2_or2_1 _16511_ (
    .A(_06561_),
    .B(_06653_),
    .X(data_o_28_)
  );
  sg13g2_o21ai_1 _16512_ (
    .A1(addr_i_2_),
    .A2(_01421_),
    .B1(_03964_),
    .Y(_06654_)
  );
  sg13g2_nand2_1 _16513_ (
    .A(addr_i_3_),
    .B(_06654_),
    .Y(_06655_)
  );
  sg13g2_o21ai_1 _16514_ (
    .A1(_07547_),
    .A2(_00626_),
    .B1(addr_i_2_),
    .Y(_06656_)
  );
  sg13g2_a21oi_1 _16515_ (
    .A1(_06655_),
    .A2(_06656_),
    .B1(addr_i_4_),
    .Y(_06657_)
  );
  sg13g2_a21oi_1 _16516_ (
    .A1(_00414_),
    .A2(_02165_),
    .B1(_00565_),
    .Y(_06658_)
  );
  sg13g2_a22oi_1 _16517_ (
    .A1(_01935_),
    .A2(_04993_),
    .B1(_06658_),
    .B2(_06010_),
    .Y(_06659_)
  );
  sg13g2_o21ai_1 _16518_ (
    .A1(_06630_),
    .A2(_06659_),
    .B1(_00458_),
    .Y(_06660_)
  );
  sg13g2_o21ai_1 _16519_ (
    .A1(_06657_),
    .A2(_06660_),
    .B1(addr_i_8_),
    .Y(_06661_)
  );
  sg13g2_nand2_1 _16520_ (
    .A(_09476_),
    .B(_05780_),
    .Y(_06663_)
  );
  sg13g2_o21ai_1 _16521_ (
    .A1(_01290_),
    .A2(_03497_),
    .B1(_08431_),
    .Y(_06664_)
  );
  sg13g2_a21o_1 _16522_ (
    .A1(_05877_),
    .A2(_06663_),
    .B1(_06664_),
    .X(_06665_)
  );
  sg13g2_a21oi_1 _16523_ (
    .A1(_00565_),
    .A2(_00328_),
    .B1(_00743_),
    .Y(_06666_)
  );
  sg13g2_a21oi_1 _16524_ (
    .A1(_03235_),
    .A2(_06666_),
    .B1(addr_i_4_),
    .Y(_06667_)
  );
  sg13g2_a22oi_1 _16525_ (
    .A1(addr_i_4_),
    .A2(_09448_),
    .B1(_06667_),
    .B2(_01082_),
    .Y(_06668_)
  );
  sg13g2_a22oi_1 _16526_ (
    .A1(_00277_),
    .A2(_06665_),
    .B1(_06668_),
    .B2(addr_i_9_),
    .Y(_06669_)
  );
  sg13g2_nand2_1 _16527_ (
    .A(_02732_),
    .B(_01580_),
    .Y(_06670_)
  );
  sg13g2_a22oi_1 _16528_ (
    .A1(_02105_),
    .A2(_02874_),
    .B1(_09459_),
    .B2(_00261_),
    .Y(_06671_)
  );
  sg13g2_a21oi_1 _16529_ (
    .A1(_00886_),
    .A2(_06670_),
    .B1(_06671_),
    .Y(_06672_)
  );
  sg13g2_a21oi_1 _16530_ (
    .A1(_03431_),
    .A2(_00531_),
    .B1(addr_i_7_),
    .Y(_06674_)
  );
  sg13g2_o21ai_1 _16531_ (
    .A1(_06672_),
    .A2(_06674_),
    .B1(addr_i_4_),
    .Y(_06675_)
  );
  sg13g2_o21ai_1 _16532_ (
    .A1(_03775_),
    .A2(_02578_),
    .B1(_04624_),
    .Y(_06676_)
  );
  sg13g2_a21oi_1 _16533_ (
    .A1(addr_i_7_),
    .A2(_06873_),
    .B1(_00595_),
    .Y(_06677_)
  );
  sg13g2_a21oi_1 _16534_ (
    .A1(addr_i_7_),
    .A2(_06676_),
    .B1(_06677_),
    .Y(_06678_)
  );
  sg13g2_nand2_1 _16535_ (
    .A(_06675_),
    .B(_06678_),
    .Y(_06679_)
  );
  sg13g2_nor3_1 _16536_ (
    .A(_01282_),
    .B(_00401_),
    .C(_00542_),
    .Y(_06680_)
  );
  sg13g2_a21oi_1 _16537_ (
    .A1(addr_i_3_),
    .A2(_03129_),
    .B1(_06680_),
    .Y(_06681_)
  );
  sg13g2_o21ai_1 _16538_ (
    .A1(_04672_),
    .A2(_06681_),
    .B1(addr_i_9_),
    .Y(_06682_)
  );
  sg13g2_a21oi_1 _16539_ (
    .A1(_01872_),
    .A2(_06324_),
    .B1(addr_i_4_),
    .Y(_06683_)
  );
  sg13g2_nor2_1 _16540_ (
    .A(_01803_),
    .B(_06683_),
    .Y(_06685_)
  );
  sg13g2_o21ai_1 _16541_ (
    .A1(_03720_),
    .A2(_05709_),
    .B1(addr_i_5_),
    .Y(_06686_)
  );
  sg13g2_a21oi_1 _16542_ (
    .A1(_06685_),
    .A2(_06686_),
    .B1(_01082_),
    .Y(_06687_)
  );
  sg13g2_a22oi_1 _16543_ (
    .A1(addr_i_8_),
    .A2(_06679_),
    .B1(_06682_),
    .B2(_06687_),
    .Y(_06688_)
  );
  sg13g2_a22oi_1 _16544_ (
    .A1(_06661_),
    .A2(_06669_),
    .B1(addr_i_10_),
    .B2(_06688_),
    .Y(_06689_)
  );
  sg13g2_nand2_1 _16545_ (
    .A(_00960_),
    .B(_07038_),
    .Y(_06690_)
  );
  sg13g2_a21o_1 _16546_ (
    .A1(_00006_),
    .A2(_09508_),
    .B1(addr_i_4_),
    .X(_06691_)
  );
  sg13g2_a21oi_1 _16547_ (
    .A1(_06690_),
    .A2(_06691_),
    .B1(addr_i_5_),
    .Y(_06692_)
  );
  sg13g2_nor2_1 _16548_ (
    .A(_01680_),
    .B(_04316_),
    .Y(_06693_)
  );
  sg13g2_nor2_1 _16549_ (
    .A(_09105_),
    .B(_06693_),
    .Y(_06694_)
  );
  sg13g2_o21ai_1 _16550_ (
    .A1(_06692_),
    .A2(_06694_),
    .B1(addr_i_2_),
    .Y(_06696_)
  );
  sg13g2_a22oi_1 _16551_ (
    .A1(addr_i_4_),
    .A2(_04572_),
    .B1(_00057_),
    .B2(addr_i_3_),
    .Y(_06697_)
  );
  sg13g2_a221oi_1 _16552_ (
    .A1(_09497_),
    .A2(_05236_),
    .B1(_01252_),
    .B2(_01228_),
    .C1(_04461_),
    .Y(_06698_)
  );
  sg13g2_nor2_1 _16553_ (
    .A(_06697_),
    .B(_06698_),
    .Y(_06699_)
  );
  sg13g2_a221oi_1 _16554_ (
    .A1(_04442_),
    .A2(_03572_),
    .B1(_06699_),
    .B2(_00146_),
    .C1(_01043_),
    .Y(_06700_)
  );
  sg13g2_nand3_1 _16555_ (
    .A(addr_i_3_),
    .B(addr_i_2_),
    .C(_07038_),
    .Y(_06701_)
  );
  sg13g2_nand3_1 _16556_ (
    .A(_04450_),
    .B(addr_i_7_),
    .C(_09371_),
    .Y(_06702_)
  );
  sg13g2_a21oi_1 _16557_ (
    .A1(_06701_),
    .A2(_06702_),
    .B1(addr_i_5_),
    .Y(_06703_)
  );
  sg13g2_a221oi_1 _16558_ (
    .A1(_06054_),
    .A2(_04572_),
    .B1(_03348_),
    .B2(_09127_),
    .C1(_06703_),
    .Y(_06704_)
  );
  sg13g2_a21oi_1 _16559_ (
    .A1(_00506_),
    .A2(_00140_),
    .B1(addr_i_7_),
    .Y(_06705_)
  );
  sg13g2_a22oi_1 _16560_ (
    .A1(_00645_),
    .A2(_06115_),
    .B1(_06705_),
    .B2(addr_i_4_),
    .Y(_06707_)
  );
  sg13g2_a21oi_1 _16561_ (
    .A1(addr_i_4_),
    .A2(_06704_),
    .B1(_06707_),
    .Y(_06708_)
  );
  sg13g2_a22oi_1 _16562_ (
    .A1(_00239_),
    .A2(_03572_),
    .B1(_06708_),
    .B2(addr_i_8_),
    .Y(_06709_)
  );
  sg13g2_a22oi_1 _16563_ (
    .A1(_06696_),
    .A2(_06700_),
    .B1(_00925_),
    .B2(_06709_),
    .Y(_06710_)
  );
  sg13g2_nand2_1 _16564_ (
    .A(_02081_),
    .B(_02807_),
    .Y(_06711_)
  );
  sg13g2_nor3_1 _16565_ (
    .A(_07270_),
    .B(_00077_),
    .C(_00279_),
    .Y(_06712_)
  );
  sg13g2_a22oi_1 _16566_ (
    .A1(_09474_),
    .A2(_06711_),
    .B1(_06712_),
    .B2(addr_i_8_),
    .Y(_06713_)
  );
  sg13g2_a21oi_1 _16567_ (
    .A1(addr_i_3_),
    .A2(_00848_),
    .B1(_01846_),
    .Y(_06714_)
  );
  sg13g2_nor2_1 _16568_ (
    .A(addr_i_6_),
    .B(_06714_),
    .Y(_06715_)
  );
  sg13g2_a21oi_1 _16569_ (
    .A1(_06070_),
    .A2(_00894_),
    .B1(_00497_),
    .Y(_06716_)
  );
  sg13g2_o21ai_1 _16570_ (
    .A1(_06715_),
    .A2(_06716_),
    .B1(addr_i_7_),
    .Y(_06719_)
  );
  sg13g2_and2_1 _16571_ (
    .A(_02529_),
    .B(_02048_),
    .X(_06720_)
  );
  sg13g2_o21ai_1 _16572_ (
    .A1(addr_i_3_),
    .A2(_06720_),
    .B1(_01921_),
    .Y(_06721_)
  );
  sg13g2_a22oi_1 _16573_ (
    .A1(_00822_),
    .A2(_06094_),
    .B1(_02226_),
    .B2(_03980_),
    .Y(_06722_)
  );
  sg13g2_o21ai_1 _16574_ (
    .A1(_00059_),
    .A2(_02103_),
    .B1(_00927_),
    .Y(_06723_)
  );
  sg13g2_a221oi_1 _16575_ (
    .A1(_01881_),
    .A2(_02598_),
    .B1(_06723_),
    .B2(addr_i_6_),
    .C1(_00112_),
    .Y(_06724_)
  );
  sg13g2_o21ai_1 _16576_ (
    .A1(addr_i_7_),
    .A2(_06722_),
    .B1(_06724_),
    .Y(_06725_)
  );
  sg13g2_a21oi_1 _16577_ (
    .A1(addr_i_7_),
    .A2(_06721_),
    .B1(_06725_),
    .Y(_06726_)
  );
  sg13g2_a22oi_1 _16578_ (
    .A1(_06713_),
    .A2(_06719_),
    .B1(_06726_),
    .B2(_06652_),
    .Y(_06727_)
  );
  sg13g2_or3_1 _16579_ (
    .A(addr_i_11_),
    .B(_06710_),
    .C(_06727_),
    .X(_06728_)
  );
  sg13g2_nor3_1 _16580_ (
    .A(_00507_),
    .B(_00770_),
    .C(_01007_),
    .Y(_06730_)
  );
  sg13g2_o21ai_1 _16581_ (
    .A1(_01645_),
    .A2(_06730_),
    .B1(_01350_),
    .Y(_06731_)
  );
  sg13g2_o21ai_1 _16582_ (
    .A1(_00820_),
    .A2(_01754_),
    .B1(_02695_),
    .Y(_06732_)
  );
  sg13g2_nand2_1 _16583_ (
    .A(addr_i_8_),
    .B(_01948_),
    .Y(_06733_)
  );
  sg13g2_o21ai_1 _16584_ (
    .A1(addr_i_7_),
    .A2(_09497_),
    .B1(addr_i_2_),
    .Y(_06734_)
  );
  sg13g2_nand2_1 _16585_ (
    .A(_00072_),
    .B(_00292_),
    .Y(_06735_)
  );
  sg13g2_a21oi_1 _16586_ (
    .A1(_06734_),
    .A2(_06735_),
    .B1(addr_i_6_),
    .Y(_06736_)
  );
  sg13g2_a22oi_1 _16587_ (
    .A1(_01475_),
    .A2(_06732_),
    .B1(_06733_),
    .B2(_06736_),
    .Y(_06737_)
  );
  sg13g2_a21oi_1 _16588_ (
    .A1(_01729_),
    .A2(_01499_),
    .B1(_02271_),
    .Y(_06738_)
  );
  sg13g2_o21ai_1 _16589_ (
    .A1(_02170_),
    .A2(_06738_),
    .B1(_01794_),
    .Y(_06739_)
  );
  sg13g2_a22oi_1 _16590_ (
    .A1(_01144_),
    .A2(_01060_),
    .B1(_00168_),
    .B2(_02297_),
    .Y(_06741_)
  );
  sg13g2_o21ai_1 _16591_ (
    .A1(_05292_),
    .A2(_02935_),
    .B1(addr_i_7_),
    .Y(_06742_)
  );
  sg13g2_nand3_1 _16592_ (
    .A(_03820_),
    .B(_03993_),
    .C(_08553_),
    .Y(_06743_)
  );
  sg13g2_a21oi_1 _16593_ (
    .A1(_06742_),
    .A2(_06743_),
    .B1(addr_i_4_),
    .Y(_06744_)
  );
  sg13g2_nor3_1 _16594_ (
    .A(addr_i_8_),
    .B(_06741_),
    .C(_06744_),
    .Y(_06745_)
  );
  sg13g2_a22oi_1 _16595_ (
    .A1(_06737_),
    .A2(_06739_),
    .B1(_06745_),
    .B2(addr_i_9_),
    .Y(_06746_)
  );
  sg13g2_and3_1 _16596_ (
    .A(addr_i_9_),
    .B(_04604_),
    .C(_01668_),
    .X(_06747_)
  );
  sg13g2_o21ai_1 _16597_ (
    .A1(_06746_),
    .A2(_06747_),
    .B1(_00511_),
    .Y(_06748_)
  );
  sg13g2_nand3_1 _16598_ (
    .A(addr_i_11_),
    .B(_06731_),
    .C(_06748_),
    .Y(_06749_)
  );
  sg13g2_o21ai_1 _16599_ (
    .A1(_06689_),
    .A2(_06728_),
    .B1(_06749_),
    .Y(_06750_)
  );
  sg13g2_nand2_1 _16600_ (
    .A(_04429_),
    .B(_01438_),
    .Y(_06752_)
  );
  sg13g2_o21ai_1 _16601_ (
    .A1(addr_i_4_),
    .A2(_08188_),
    .B1(addr_i_3_),
    .Y(_06753_)
  );
  sg13g2_a21oi_1 _16602_ (
    .A1(_04451_),
    .A2(_06753_),
    .B1(addr_i_2_),
    .Y(_06754_)
  );
  sg13g2_a21oi_1 _16603_ (
    .A1(_01336_),
    .A2(_06752_),
    .B1(_06754_),
    .Y(_06755_)
  );
  sg13g2_o21ai_1 _16604_ (
    .A1(addr_i_3_),
    .A2(_09504_),
    .B1(_01967_),
    .Y(_06756_)
  );
  sg13g2_a221oi_1 _16605_ (
    .A1(_00157_),
    .A2(_00096_),
    .B1(_06756_),
    .B2(addr_i_2_),
    .C1(addr_i_5_),
    .Y(_06757_)
  );
  sg13g2_a21oi_1 _16606_ (
    .A1(addr_i_5_),
    .A2(_06755_),
    .B1(_06757_),
    .Y(_06758_)
  );
  sg13g2_o21ai_1 _16607_ (
    .A1(_09205_),
    .A2(_06983_),
    .B1(_00677_),
    .Y(_06759_)
  );
  sg13g2_nand2_1 _16608_ (
    .A(_00763_),
    .B(_00975_),
    .Y(_06760_)
  );
  sg13g2_nor3_1 _16609_ (
    .A(addr_i_4_),
    .B(addr_i_5_),
    .C(_00086_),
    .Y(_06761_)
  );
  sg13g2_o21ai_1 _16610_ (
    .A1(_06760_),
    .A2(_06761_),
    .B1(_00091_),
    .Y(_06763_)
  );
  sg13g2_o21ai_1 _16611_ (
    .A1(_00573_),
    .A2(_04016_),
    .B1(_06763_),
    .Y(_06764_)
  );
  sg13g2_o21ai_1 _16612_ (
    .A1(_03358_),
    .A2(_00533_),
    .B1(_05427_),
    .Y(_06765_)
  );
  sg13g2_a221oi_1 _16613_ (
    .A1(addr_i_2_),
    .A2(_06759_),
    .B1(_06764_),
    .B2(_03260_),
    .C1(_06765_),
    .Y(_06766_)
  );
  sg13g2_nor2_1 _16614_ (
    .A(addr_i_8_),
    .B(_06766_),
    .Y(_06767_)
  );
  sg13g2_a22oi_1 _16615_ (
    .A1(addr_i_8_),
    .A2(_06758_),
    .B1(_06767_),
    .B2(_02221_),
    .Y(_06768_)
  );
  sg13g2_o21ai_1 _16616_ (
    .A1(addr_i_2_),
    .A2(_04747_),
    .B1(_06895_),
    .Y(_06769_)
  );
  sg13g2_nand2_1 _16617_ (
    .A(_01861_),
    .B(_00943_),
    .Y(_06770_)
  );
  sg13g2_a21oi_1 _16618_ (
    .A1(_07724_),
    .A2(_06339_),
    .B1(_03292_),
    .Y(_06771_)
  );
  sg13g2_a22oi_1 _16619_ (
    .A1(_00061_),
    .A2(_06769_),
    .B1(_06770_),
    .B2(_06771_),
    .Y(_06772_)
  );
  sg13g2_nand2_1 _16620_ (
    .A(_01729_),
    .B(_01060_),
    .Y(_06774_)
  );
  sg13g2_nand3_1 _16621_ (
    .A(addr_i_6_),
    .B(_00692_),
    .C(_01872_),
    .Y(_06775_)
  );
  sg13g2_a21oi_1 _16622_ (
    .A1(_09478_),
    .A2(_06775_),
    .B1(addr_i_4_),
    .Y(_06776_)
  );
  sg13g2_a22oi_1 _16623_ (
    .A1(addr_i_4_),
    .A2(_06774_),
    .B1(_06776_),
    .B2(_06497_),
    .Y(_06777_)
  );
  sg13g2_nor2_1 _16624_ (
    .A(_01391_),
    .B(_06777_),
    .Y(_06778_)
  );
  sg13g2_nand2_1 _16625_ (
    .A(_07812_),
    .B(_03172_),
    .Y(_06779_)
  );
  sg13g2_nand3_1 _16626_ (
    .A(_04162_),
    .B(_06779_),
    .C(_06528_),
    .Y(_06780_)
  );
  sg13g2_a22oi_1 _16627_ (
    .A1(addr_i_4_),
    .A2(_06780_),
    .B1(_03070_),
    .B2(_00474_),
    .Y(_06781_)
  );
  sg13g2_nor2_1 _16628_ (
    .A(addr_i_7_),
    .B(_06781_),
    .Y(_06782_)
  );
  sg13g2_a21oi_1 _16629_ (
    .A1(_03226_),
    .A2(_05775_),
    .B1(_03930_),
    .Y(_06783_)
  );
  sg13g2_a22oi_1 _16630_ (
    .A1(_00073_),
    .A2(_02119_),
    .B1(_06783_),
    .B2(_00779_),
    .Y(_06785_)
  );
  sg13g2_nor3_1 _16631_ (
    .A(addr_i_8_),
    .B(_06782_),
    .C(_06785_),
    .Y(_06786_)
  );
  sg13g2_nor4_1 _16632_ (
    .A(_01211_),
    .B(_06772_),
    .C(_06778_),
    .D(_06786_),
    .Y(_06787_)
  );
  sg13g2_nor3_1 _16633_ (
    .A(addr_i_11_),
    .B(_06768_),
    .C(_06787_),
    .Y(_06788_)
  );
  sg13g2_nand2_1 _16634_ (
    .A(_03575_),
    .B(_00353_),
    .Y(_06789_)
  );
  sg13g2_nand2_1 _16635_ (
    .A(_03908_),
    .B(_04793_),
    .Y(_06790_)
  );
  sg13g2_nor2_1 _16636_ (
    .A(addr_i_3_),
    .B(_09448_),
    .Y(_06791_)
  );
  sg13g2_a22oi_1 _16637_ (
    .A1(addr_i_3_),
    .A2(_06790_),
    .B1(_06791_),
    .B2(_00360_),
    .Y(_06792_)
  );
  sg13g2_a22oi_1 _16638_ (
    .A1(_01240_),
    .A2(_06789_),
    .B1(_06792_),
    .B2(addr_i_8_),
    .Y(_06793_)
  );
  sg13g2_nand3_1 _16639_ (
    .A(addr_i_3_),
    .B(_02898_),
    .C(_00878_),
    .Y(_06794_)
  );
  sg13g2_nand3_1 _16640_ (
    .A(_05867_),
    .B(_01290_),
    .C(_01029_),
    .Y(_06796_)
  );
  sg13g2_a221oi_1 _16641_ (
    .A1(_04052_),
    .A2(_02410_),
    .B1(_06794_),
    .B2(_06796_),
    .C1(_00629_),
    .Y(_06797_)
  );
  sg13g2_nor2_1 _16642_ (
    .A(_06793_),
    .B(_06797_),
    .Y(_06798_)
  );
  sg13g2_nand3_1 _16643_ (
    .A(_06895_),
    .B(_02810_),
    .C(_05012_),
    .Y(_06799_)
  );
  sg13g2_a21oi_1 _16644_ (
    .A1(_01367_),
    .A2(_00430_),
    .B1(addr_i_5_),
    .Y(_06800_)
  );
  sg13g2_a21oi_1 _16645_ (
    .A1(addr_i_3_),
    .A2(_06799_),
    .B1(_06800_),
    .Y(_06801_)
  );
  sg13g2_nor2_1 _16646_ (
    .A(_01082_),
    .B(_06801_),
    .Y(_06802_)
  );
  sg13g2_a21oi_1 _16647_ (
    .A1(_03431_),
    .A2(_01709_),
    .B1(_08399_),
    .Y(_06803_)
  );
  sg13g2_a21oi_1 _16648_ (
    .A1(addr_i_4_),
    .A2(_06884_),
    .B1(addr_i_3_),
    .Y(_06804_)
  );
  sg13g2_a22oi_1 _16649_ (
    .A1(_01500_),
    .A2(_03497_),
    .B1(_02542_),
    .B2(_06804_),
    .Y(_06805_)
  );
  sg13g2_nand2_1 _16650_ (
    .A(_01118_),
    .B(_06805_),
    .Y(_06807_)
  );
  sg13g2_o21ai_1 _16651_ (
    .A1(_06803_),
    .A2(_06807_),
    .B1(addr_i_9_),
    .Y(_06808_)
  );
  sg13g2_a22oi_1 _16652_ (
    .A1(addr_i_7_),
    .A2(_06798_),
    .B1(_06802_),
    .B2(_06808_),
    .Y(_06809_)
  );
  sg13g2_a21oi_1 _16653_ (
    .A1(_00391_),
    .A2(_03845_),
    .B1(_01234_),
    .Y(_06810_)
  );
  sg13g2_o21ai_1 _16654_ (
    .A1(_02935_),
    .A2(_06033_),
    .B1(addr_i_4_),
    .Y(_06811_)
  );
  sg13g2_a21oi_1 _16655_ (
    .A1(_00545_),
    .A2(_06811_),
    .B1(_00825_),
    .Y(_06812_)
  );
  sg13g2_a21oi_1 _16656_ (
    .A1(_01103_),
    .A2(_02708_),
    .B1(_01125_),
    .Y(_06813_)
  );
  sg13g2_a21oi_1 _16657_ (
    .A1(_03993_),
    .A2(_03243_),
    .B1(_06813_),
    .Y(_06814_)
  );
  sg13g2_nor2_1 _16658_ (
    .A(addr_i_7_),
    .B(_06814_),
    .Y(_06815_)
  );
  sg13g2_nor4_1 _16659_ (
    .A(_00214_),
    .B(_06810_),
    .C(_06812_),
    .D(_06815_),
    .Y(_06816_)
  );
  sg13g2_nor2_1 _16660_ (
    .A(addr_i_3_),
    .B(_05425_),
    .Y(_06818_)
  );
  sg13g2_o21ai_1 _16661_ (
    .A1(_00850_),
    .A2(_06818_),
    .B1(_00169_),
    .Y(_06819_)
  );
  sg13g2_nand2_1 _16662_ (
    .A(_00845_),
    .B(_02807_),
    .Y(_06820_)
  );
  sg13g2_a22oi_1 _16663_ (
    .A1(_00529_),
    .A2(_06820_),
    .B1(_04791_),
    .B2(addr_i_9_),
    .Y(_06821_)
  );
  sg13g2_a21oi_1 _16664_ (
    .A1(_06032_),
    .A2(_01029_),
    .B1(_00700_),
    .Y(_06822_)
  );
  sg13g2_o21ai_1 _16665_ (
    .A1(_01803_),
    .A2(_06822_),
    .B1(_08708_),
    .Y(_06823_)
  );
  sg13g2_o21ai_1 _16666_ (
    .A1(_00227_),
    .A2(_07503_),
    .B1(addr_i_6_),
    .Y(_06824_)
  );
  sg13g2_a21o_1 _16667_ (
    .A1(_06823_),
    .A2(_06824_),
    .B1(addr_i_7_),
    .X(_06825_)
  );
  sg13g2_nand3_1 _16668_ (
    .A(_06819_),
    .B(_06821_),
    .C(_06825_),
    .Y(_06826_)
  );
  sg13g2_nand2b_1 _16669_ (
    .A_N(_06816_),
    .B(_06826_),
    .Y(_06827_)
  );
  sg13g2_o21ai_1 _16670_ (
    .A1(_06809_),
    .A2(_06827_),
    .B1(_01774_),
    .Y(_06830_)
  );
  sg13g2_nand2_1 _16671_ (
    .A(_02732_),
    .B(_01588_),
    .Y(_06831_)
  );
  sg13g2_a21oi_1 _16672_ (
    .A1(_04451_),
    .A2(_02895_),
    .B1(addr_i_2_),
    .Y(_06832_)
  );
  sg13g2_a22oi_1 _16673_ (
    .A1(_07824_),
    .A2(_06831_),
    .B1(_06832_),
    .B2(_00206_),
    .Y(_06833_)
  );
  sg13g2_nand2_1 _16674_ (
    .A(_00884_),
    .B(_01749_),
    .Y(_06834_)
  );
  sg13g2_o21ai_1 _16675_ (
    .A1(_03809_),
    .A2(_02196_),
    .B1(addr_i_4_),
    .Y(_06835_)
  );
  sg13g2_a221oi_1 _16676_ (
    .A1(addr_i_3_),
    .A2(_00441_),
    .B1(_06835_),
    .B2(_00445_),
    .C1(addr_i_6_),
    .Y(_06836_)
  );
  sg13g2_a22oi_1 _16677_ (
    .A1(_05600_),
    .A2(_06834_),
    .B1(_06836_),
    .B2(addr_i_8_),
    .Y(_06837_)
  );
  sg13g2_o21ai_1 _16678_ (
    .A1(_01475_),
    .A2(_06833_),
    .B1(_06837_),
    .Y(_06838_)
  );
  sg13g2_nor2_1 _16679_ (
    .A(_00768_),
    .B(_00718_),
    .Y(_06839_)
  );
  sg13g2_o21ai_1 _16680_ (
    .A1(_05195_),
    .A2(_06839_),
    .B1(_05236_),
    .Y(_06841_)
  );
  sg13g2_o21ai_1 _16681_ (
    .A1(_02569_),
    .A2(_06179_),
    .B1(_06841_),
    .Y(_06842_)
  );
  sg13g2_o21ai_1 _16682_ (
    .A1(addr_i_3_),
    .A2(_03233_),
    .B1(_01709_),
    .Y(_06843_)
  );
  sg13g2_a21oi_1 _16683_ (
    .A1(_07326_),
    .A2(_00863_),
    .B1(_02387_),
    .Y(_06844_)
  );
  sg13g2_o21ai_1 _16684_ (
    .A1(_00252_),
    .A2(_01943_),
    .B1(_06364_),
    .Y(_06845_)
  );
  sg13g2_nand3_1 _16685_ (
    .A(addr_i_7_),
    .B(_00704_),
    .C(_06845_),
    .Y(_06846_)
  );
  sg13g2_a22oi_1 _16686_ (
    .A1(addr_i_4_),
    .A2(_06843_),
    .B1(_06844_),
    .B2(_06846_),
    .Y(_06847_)
  );
  sg13g2_nor3_1 _16687_ (
    .A(_01559_),
    .B(_06842_),
    .C(_06847_),
    .Y(_06848_)
  );
  sg13g2_nor2_1 _16688_ (
    .A(_09315_),
    .B(_06848_),
    .Y(_06849_)
  );
  sg13g2_o21ai_1 _16689_ (
    .A1(_06419_),
    .A2(_05318_),
    .B1(_00940_),
    .Y(_06850_)
  );
  sg13g2_a21oi_1 _16690_ (
    .A1(_01339_),
    .A2(_00687_),
    .B1(_02577_),
    .Y(_06852_)
  );
  sg13g2_nand3_1 _16691_ (
    .A(_04494_),
    .B(_09371_),
    .C(_00926_),
    .Y(_06853_)
  );
  sg13g2_o21ai_1 _16692_ (
    .A1(_00406_),
    .A2(_00961_),
    .B1(_00025_),
    .Y(_06854_)
  );
  sg13g2_a22oi_1 _16693_ (
    .A1(addr_i_3_),
    .A2(_06853_),
    .B1(_06854_),
    .B2(_04681_),
    .Y(_06855_)
  );
  sg13g2_nor2_1 _16694_ (
    .A(addr_i_5_),
    .B(_06855_),
    .Y(_06856_)
  );
  sg13g2_a22oi_1 _16695_ (
    .A1(addr_i_7_),
    .A2(_06850_),
    .B1(_06852_),
    .B2(_06856_),
    .Y(_06857_)
  );
  sg13g2_o21ai_1 _16696_ (
    .A1(_01507_),
    .A2(_02623_),
    .B1(addr_i_4_),
    .Y(_06858_)
  );
  sg13g2_nand2_1 _16697_ (
    .A(_00249_),
    .B(_06858_),
    .Y(_06859_)
  );
  sg13g2_nor2_1 _16698_ (
    .A(_01659_),
    .B(_01746_),
    .Y(_06860_)
  );
  sg13g2_o21ai_1 _16699_ (
    .A1(_00127_),
    .A2(_01782_),
    .B1(_05070_),
    .Y(_06861_)
  );
  sg13g2_a21oi_1 _16700_ (
    .A1(_06860_),
    .A2(_06861_),
    .B1(addr_i_6_),
    .Y(_06863_)
  );
  sg13g2_a22oi_1 _16701_ (
    .A1(_01480_),
    .A2(_06859_),
    .B1(_06863_),
    .B2(addr_i_8_),
    .Y(_06864_)
  );
  sg13g2_a22oi_1 _16702_ (
    .A1(addr_i_8_),
    .A2(_06857_),
    .B1(_06864_),
    .B2(addr_i_9_),
    .Y(_06865_)
  );
  sg13g2_a21o_1 _16703_ (
    .A1(_06838_),
    .A2(_06849_),
    .B1(_06865_),
    .X(_06866_)
  );
  sg13g2_a21oi_1 _16704_ (
    .A1(_01277_),
    .A2(_00844_),
    .B1(_05512_),
    .Y(_06867_)
  );
  sg13g2_o21ai_1 _16705_ (
    .A1(_07149_),
    .A2(_06867_),
    .B1(_03771_),
    .Y(_06868_)
  );
  sg13g2_o21ai_1 _16706_ (
    .A1(_01202_),
    .A2(_06839_),
    .B1(addr_i_6_),
    .Y(_06869_)
  );
  sg13g2_o21ai_1 _16707_ (
    .A1(_00617_),
    .A2(_00945_),
    .B1(addr_i_3_),
    .Y(_06870_)
  );
  sg13g2_a21oi_1 _16708_ (
    .A1(_06869_),
    .A2(_06870_),
    .B1(_07614_),
    .Y(_06871_)
  );
  sg13g2_a21oi_1 _16709_ (
    .A1(_01861_),
    .A2(_06868_),
    .B1(_06871_),
    .Y(_06872_)
  );
  sg13g2_or3_1 _16710_ (
    .A(addr_i_3_),
    .B(_01779_),
    .C(_09094_),
    .X(_06874_)
  );
  sg13g2_nor2_1 _16711_ (
    .A(_02949_),
    .B(_04139_),
    .Y(_06875_)
  );
  sg13g2_a21oi_1 _16712_ (
    .A1(addr_i_3_),
    .A2(_06875_),
    .B1(_08830_),
    .Y(_06876_)
  );
  sg13g2_a21oi_1 _16713_ (
    .A1(addr_i_5_),
    .A2(_05910_),
    .B1(_05324_),
    .Y(_06877_)
  );
  sg13g2_o21ai_1 _16714_ (
    .A1(_00205_),
    .A2(_06877_),
    .B1(addr_i_2_),
    .Y(_06878_)
  );
  sg13g2_a21oi_1 _16715_ (
    .A1(_04916_),
    .A2(_06878_),
    .B1(_07403_),
    .Y(_06879_)
  );
  sg13g2_a22oi_1 _16716_ (
    .A1(_06874_),
    .A2(_06876_),
    .B1(addr_i_9_),
    .B2(_06879_),
    .Y(_06880_)
  );
  sg13g2_nor3_1 _16717_ (
    .A(addr_i_2_),
    .B(_00006_),
    .C(_01208_),
    .Y(_06881_)
  );
  sg13g2_nand2_1 _16718_ (
    .A(_00764_),
    .B(_03350_),
    .Y(_06882_)
  );
  sg13g2_nor4_1 _16719_ (
    .A(_02598_),
    .B(_03742_),
    .C(_06881_),
    .D(_06882_),
    .Y(_06883_)
  );
  sg13g2_a22oi_1 _16720_ (
    .A1(_00702_),
    .A2(_01795_),
    .B1(_00343_),
    .B2(addr_i_7_),
    .Y(_06885_)
  );
  sg13g2_o21ai_1 _16721_ (
    .A1(_09513_),
    .A2(_04475_),
    .B1(_05648_),
    .Y(_06886_)
  );
  sg13g2_nor2_1 _16722_ (
    .A(_06885_),
    .B(_06886_),
    .Y(_06887_)
  );
  sg13g2_o21ai_1 _16723_ (
    .A1(addr_i_4_),
    .A2(_06883_),
    .B1(_06887_),
    .Y(_06888_)
  );
  sg13g2_o21ai_1 _16724_ (
    .A1(_00998_),
    .A2(_06877_),
    .B1(addr_i_2_),
    .Y(_06889_)
  );
  sg13g2_nand4_1 _16725_ (
    .A(_02708_),
    .B(_03324_),
    .C(_03745_),
    .D(_06889_),
    .Y(_06890_)
  );
  sg13g2_o21ai_1 _16726_ (
    .A1(_01070_),
    .A2(_02191_),
    .B1(_01301_),
    .Y(_06891_)
  );
  sg13g2_nor2_1 _16727_ (
    .A(addr_i_6_),
    .B(_00384_),
    .Y(_06892_)
  );
  sg13g2_o21ai_1 _16728_ (
    .A1(_01182_),
    .A2(_06892_),
    .B1(addr_i_8_),
    .Y(_06893_)
  );
  sg13g2_o21ai_1 _16729_ (
    .A1(addr_i_4_),
    .A2(_01580_),
    .B1(_08410_),
    .Y(_06894_)
  );
  sg13g2_nand2b_1 _16730_ (
    .A_N(_06893_),
    .B(_06894_),
    .Y(_06896_)
  );
  sg13g2_a221oi_1 _16731_ (
    .A1(_05822_),
    .A2(_06890_),
    .B1(_06891_),
    .B2(_07149_),
    .C1(_06896_),
    .Y(_06897_)
  );
  sg13g2_a22oi_1 _16732_ (
    .A1(_07293_),
    .A2(_06888_),
    .B1(_06897_),
    .B2(_01351_),
    .Y(_06898_)
  );
  sg13g2_a22oi_1 _16733_ (
    .A1(_06872_),
    .A2(_06880_),
    .B1(_06898_),
    .B2(addr_i_10_),
    .Y(_06899_)
  );
  sg13g2_a21o_1 _16734_ (
    .A1(addr_i_10_),
    .A2(_06866_),
    .B1(_06899_),
    .X(_06900_)
  );
  sg13g2_a221oi_1 _16735_ (
    .A1(_06788_),
    .A2(_06830_),
    .B1(_06900_),
    .B2(addr_i_11_),
    .C1(addr_i_12_),
    .Y(_06901_)
  );
  sg13g2_a21oi_1 _16736_ (
    .A1(addr_i_12_),
    .A2(_06750_),
    .B1(_06901_),
    .Y(data_o_29_)
  );
  sg13g2_a22oi_1 _16737_ (
    .A1(_02297_),
    .A2(_03348_),
    .B1(_02380_),
    .B2(_02759_),
    .Y(_06902_)
  );
  sg13g2_a21oi_1 _16738_ (
    .A1(_01252_),
    .A2(_02920_),
    .B1(addr_i_3_),
    .Y(_06903_)
  );
  sg13g2_a21oi_1 _16739_ (
    .A1(_09510_),
    .A2(_01709_),
    .B1(_08388_),
    .Y(_06904_)
  );
  sg13g2_nor4_1 _16740_ (
    .A(addr_i_7_),
    .B(_00268_),
    .C(_06903_),
    .D(_06904_),
    .Y(_06906_)
  );
  sg13g2_nor3_1 _16741_ (
    .A(_00548_),
    .B(_01986_),
    .C(_04939_),
    .Y(_06907_)
  );
  sg13g2_nor4_1 _16742_ (
    .A(addr_i_8_),
    .B(_06902_),
    .C(_06906_),
    .D(_06907_),
    .Y(_06908_)
  );
  sg13g2_nand2_1 _16743_ (
    .A(_04162_),
    .B(_00442_),
    .Y(_06909_)
  );
  sg13g2_nand2b_1 _16744_ (
    .A_N(_00854_),
    .B(_06909_),
    .Y(_06910_)
  );
  sg13g2_a221oi_1 _16745_ (
    .A1(addr_i_2_),
    .A2(_05081_),
    .B1(_05739_),
    .B2(addr_i_3_),
    .C1(_01517_),
    .Y(_06911_)
  );
  sg13g2_o21ai_1 _16746_ (
    .A1(_00901_),
    .A2(_06261_),
    .B1(addr_i_4_),
    .Y(_06912_)
  );
  sg13g2_nor2_1 _16747_ (
    .A(_00744_),
    .B(_04119_),
    .Y(_06913_)
  );
  sg13g2_o21ai_1 _16748_ (
    .A1(_06913_),
    .A2(_00279_),
    .B1(_09473_),
    .Y(_06914_)
  );
  sg13g2_nand2_1 _16749_ (
    .A(addr_i_8_),
    .B(_06914_),
    .Y(_06915_)
  );
  sg13g2_a221oi_1 _16750_ (
    .A1(_00402_),
    .A2(_06910_),
    .B1(_06911_),
    .B2(_06912_),
    .C1(_06915_),
    .Y(_06917_)
  );
  sg13g2_nor2_1 _16751_ (
    .A(_06908_),
    .B(_06917_),
    .Y(_06918_)
  );
  sg13g2_o21ai_1 _16752_ (
    .A1(addr_i_5_),
    .A2(_00605_),
    .B1(addr_i_4_),
    .Y(_06919_)
  );
  sg13g2_o21ai_1 _16753_ (
    .A1(addr_i_3_),
    .A2(_02388_),
    .B1(_06919_),
    .Y(_06920_)
  );
  sg13g2_a21oi_1 _16754_ (
    .A1(_00566_),
    .A2(_08464_),
    .B1(_00554_),
    .Y(_06921_)
  );
  sg13g2_a21o_1 _16755_ (
    .A1(_00122_),
    .A2(_06920_),
    .B1(_06921_),
    .X(_06922_)
  );
  sg13g2_o21ai_1 _16756_ (
    .A1(_01881_),
    .A2(_01759_),
    .B1(_01878_),
    .Y(_06923_)
  );
  sg13g2_nand3_1 _16757_ (
    .A(_09486_),
    .B(_02470_),
    .C(_04969_),
    .Y(_06924_)
  );
  sg13g2_nand2_1 _16758_ (
    .A(_06923_),
    .B(_06924_),
    .Y(_06925_)
  );
  sg13g2_a22oi_1 _16759_ (
    .A1(addr_i_7_),
    .A2(_06922_),
    .B1(_06925_),
    .B2(addr_i_8_),
    .Y(_06926_)
  );
  sg13g2_o21ai_1 _16760_ (
    .A1(_06795_),
    .A2(_03455_),
    .B1(addr_i_3_),
    .Y(_06928_)
  );
  sg13g2_o21ai_1 _16761_ (
    .A1(_00972_),
    .A2(_01749_),
    .B1(_06928_),
    .Y(_06929_)
  );
  sg13g2_nand2_1 _16762_ (
    .A(_00463_),
    .B(_05651_),
    .Y(_06930_)
  );
  sg13g2_a21oi_1 _16763_ (
    .A1(_00863_),
    .A2(_06930_),
    .B1(addr_i_2_),
    .Y(_06931_)
  );
  sg13g2_a22oi_1 _16764_ (
    .A1(addr_i_3_),
    .A2(_01167_),
    .B1(_06931_),
    .B2(_00416_),
    .Y(_06932_)
  );
  sg13g2_nor2_1 _16765_ (
    .A(addr_i_7_),
    .B(_06932_),
    .Y(_06933_)
  );
  sg13g2_nand3_1 _16766_ (
    .A(_09061_),
    .B(_01473_),
    .C(_03445_),
    .Y(_06934_)
  );
  sg13g2_o21ai_1 _16767_ (
    .A1(_05038_),
    .A2(_06934_),
    .B1(addr_i_8_),
    .Y(_06935_)
  );
  sg13g2_a22oi_1 _16768_ (
    .A1(_00169_),
    .A2(_06929_),
    .B1(_06933_),
    .B2(_06935_),
    .Y(_06936_)
  );
  sg13g2_nor2_1 _16769_ (
    .A(_06926_),
    .B(_06936_),
    .Y(_06937_)
  );
  sg13g2_a21oi_1 _16770_ (
    .A1(_00183_),
    .A2(_06099_),
    .B1(_09127_),
    .Y(_06940_)
  );
  sg13g2_o21ai_1 _16771_ (
    .A1(addr_i_7_),
    .A2(_07458_),
    .B1(_09226_),
    .Y(_06941_)
  );
  sg13g2_o21ai_1 _16772_ (
    .A1(addr_i_3_),
    .A2(_06940_),
    .B1(_06941_),
    .Y(_06942_)
  );
  sg13g2_nand2_1 _16773_ (
    .A(_00644_),
    .B(_01495_),
    .Y(_06943_)
  );
  sg13g2_a22oi_1 _16774_ (
    .A1(_00145_),
    .A2(_02213_),
    .B1(_01064_),
    .B2(addr_i_3_),
    .Y(_06944_)
  );
  sg13g2_a22oi_1 _16775_ (
    .A1(addr_i_3_),
    .A2(_06943_),
    .B1(_06944_),
    .B2(addr_i_4_),
    .Y(_06945_)
  );
  sg13g2_a22oi_1 _16776_ (
    .A1(addr_i_2_),
    .A2(_06942_),
    .B1(_06945_),
    .B2(_02069_),
    .Y(_06946_)
  );
  sg13g2_nor2_1 _16777_ (
    .A(_01585_),
    .B(_00946_),
    .Y(_06947_)
  );
  sg13g2_nor3_1 _16778_ (
    .A(addr_i_4_),
    .B(_00100_),
    .C(_09507_),
    .Y(_06948_)
  );
  sg13g2_a22oi_1 _16779_ (
    .A1(addr_i_4_),
    .A2(_06947_),
    .B1(_06948_),
    .B2(addr_i_3_),
    .Y(_06949_)
  );
  sg13g2_nand2_1 _16780_ (
    .A(_01438_),
    .B(_01337_),
    .Y(_06951_)
  );
  sg13g2_a22oi_1 _16781_ (
    .A1(addr_i_3_),
    .A2(_06951_),
    .B1(_02154_),
    .B2(_00119_),
    .Y(_06952_)
  );
  sg13g2_a21oi_1 _16782_ (
    .A1(_00375_),
    .A2(_05231_),
    .B1(_02420_),
    .Y(_06953_)
  );
  sg13g2_o21ai_1 _16783_ (
    .A1(addr_i_2_),
    .A2(_06952_),
    .B1(_06953_),
    .Y(_06954_)
  );
  sg13g2_o21ai_1 _16784_ (
    .A1(_06949_),
    .A2(_06954_),
    .B1(addr_i_8_),
    .Y(_06955_)
  );
  sg13g2_o21ai_1 _16785_ (
    .A1(addr_i_8_),
    .A2(_06946_),
    .B1(_06955_),
    .Y(_06956_)
  );
  sg13g2_a221oi_1 _16786_ (
    .A1(_06054_),
    .A2(_00716_),
    .B1(_02943_),
    .B2(addr_i_3_),
    .C1(_09083_),
    .Y(_06957_)
  );
  sg13g2_nand2b_1 _16787_ (
    .A_N(_09215_),
    .B(_01309_),
    .Y(_06958_)
  );
  sg13g2_a21oi_1 _16788_ (
    .A1(_01834_),
    .A2(_00819_),
    .B1(_00021_),
    .Y(_06959_)
  );
  sg13g2_nand2_1 _16789_ (
    .A(_00581_),
    .B(_07492_),
    .Y(_06960_)
  );
  sg13g2_a21oi_1 _16790_ (
    .A1(_03179_),
    .A2(_06960_),
    .B1(_00052_),
    .Y(_06962_)
  );
  sg13g2_a22oi_1 _16791_ (
    .A1(_09473_),
    .A2(_06958_),
    .B1(_06959_),
    .B2(_06962_),
    .Y(_06963_)
  );
  sg13g2_o21ai_1 _16792_ (
    .A1(_00548_),
    .A2(_06957_),
    .B1(_06963_),
    .Y(_06964_)
  );
  sg13g2_inv_1 _16793_ (
    .A(_06964_),
    .Y(_06965_)
  );
  sg13g2_a21oi_1 _16794_ (
    .A1(_00137_),
    .A2(_09477_),
    .B1(addr_i_4_),
    .Y(_06966_)
  );
  sg13g2_nor2_1 _16795_ (
    .A(_07193_),
    .B(_01659_),
    .Y(_06967_)
  );
  sg13g2_o21ai_1 _16796_ (
    .A1(addr_i_3_),
    .A2(_06967_),
    .B1(_05648_),
    .Y(_06968_)
  );
  sg13g2_o21ai_1 _16797_ (
    .A1(_06966_),
    .A2(_06968_),
    .B1(_04068_),
    .Y(_06969_)
  );
  sg13g2_o21ai_1 _16798_ (
    .A1(_01202_),
    .A2(_02923_),
    .B1(_00428_),
    .Y(_06970_)
  );
  sg13g2_or2_1 _16799_ (
    .A(_02238_),
    .B(_02847_),
    .X(_06971_)
  );
  sg13g2_a21oi_1 _16800_ (
    .A1(_02656_),
    .A2(_00832_),
    .B1(addr_i_5_),
    .Y(_06973_)
  );
  sg13g2_a22oi_1 _16801_ (
    .A1(addr_i_4_),
    .A2(_06971_),
    .B1(_06973_),
    .B2(_01711_),
    .Y(_06974_)
  );
  sg13g2_or2_1 _16802_ (
    .A(addr_i_6_),
    .B(_06974_),
    .X(_06975_)
  );
  sg13g2_and4_1 _16803_ (
    .A(_01559_),
    .B(_06969_),
    .C(_06970_),
    .D(_06975_),
    .X(_06976_)
  );
  sg13g2_a21oi_1 _16804_ (
    .A1(addr_i_8_),
    .A2(_06965_),
    .B1(_06976_),
    .Y(_06977_)
  );
  sg13g2_mux4_1 _16805_ (
    .A0(_06918_),
    .A1(_06937_),
    .A2(_06956_),
    .A3(_06977_),
    .S0(_01773_),
    .S1(_00397_),
    .X(_06978_)
  );
  sg13g2_nor2_1 _16806_ (
    .A(_00513_),
    .B(_06978_),
    .Y(_06979_)
  );
  sg13g2_nor2_1 _16807_ (
    .A(addr_i_3_),
    .B(_04658_),
    .Y(_06980_)
  );
  sg13g2_a22oi_1 _16808_ (
    .A1(_04442_),
    .A2(_04655_),
    .B1(_06980_),
    .B2(_03062_),
    .Y(_06981_)
  );
  sg13g2_o21ai_1 _16809_ (
    .A1(_00015_),
    .A2(_00503_),
    .B1(addr_i_4_),
    .Y(_06982_)
  );
  sg13g2_o21ai_1 _16810_ (
    .A1(_00190_),
    .A2(_01495_),
    .B1(_02528_),
    .Y(_06984_)
  );
  sg13g2_o21ai_1 _16811_ (
    .A1(addr_i_3_),
    .A2(_02623_),
    .B1(_03953_),
    .Y(_06985_)
  );
  sg13g2_nand2_1 _16812_ (
    .A(addr_i_2_),
    .B(_06985_),
    .Y(_06986_)
  );
  sg13g2_a21oi_1 _16813_ (
    .A1(_01504_),
    .A2(_06986_),
    .B1(addr_i_4_),
    .Y(_06987_)
  );
  sg13g2_o21ai_1 _16814_ (
    .A1(_02619_),
    .A2(_02977_),
    .B1(addr_i_3_),
    .Y(_06988_)
  );
  sg13g2_a21oi_1 _16815_ (
    .A1(_05083_),
    .A2(_06988_),
    .B1(_00497_),
    .Y(_06989_)
  );
  sg13g2_a22oi_1 _16816_ (
    .A1(_00617_),
    .A2(_06984_),
    .B1(_06987_),
    .B2(_06989_),
    .Y(_06990_)
  );
  sg13g2_nor2_1 _16817_ (
    .A(_01151_),
    .B(_06990_),
    .Y(_06991_)
  );
  sg13g2_o21ai_1 _16818_ (
    .A1(_00047_),
    .A2(_06806_),
    .B1(_03226_),
    .Y(_06992_)
  );
  sg13g2_o21ai_1 _16819_ (
    .A1(_01514_),
    .A2(_03401_),
    .B1(_01633_),
    .Y(_06993_)
  );
  sg13g2_a221oi_1 _16820_ (
    .A1(addr_i_4_),
    .A2(_02533_),
    .B1(_06992_),
    .B2(_00123_),
    .C1(_06993_),
    .Y(_06995_)
  );
  sg13g2_a22oi_1 _16821_ (
    .A1(_06981_),
    .A2(_06982_),
    .B1(_06991_),
    .B2(_06995_),
    .Y(_06996_)
  );
  sg13g2_o21ai_1 _16822_ (
    .A1(_00428_),
    .A2(_00298_),
    .B1(addr_i_5_),
    .Y(_06997_)
  );
  sg13g2_o21ai_1 _16823_ (
    .A1(_00294_),
    .A2(_09226_),
    .B1(addr_i_4_),
    .Y(_06998_)
  );
  sg13g2_a21oi_1 _16824_ (
    .A1(_06997_),
    .A2(_06998_),
    .B1(addr_i_3_),
    .Y(_06999_)
  );
  sg13g2_nand2_1 _16825_ (
    .A(_02471_),
    .B(_01672_),
    .Y(_07000_)
  );
  sg13g2_nor2_1 _16826_ (
    .A(addr_i_3_),
    .B(_04429_),
    .Y(_07001_)
  );
  sg13g2_a22oi_1 _16827_ (
    .A1(addr_i_3_),
    .A2(_07000_),
    .B1(_07001_),
    .B2(_05833_),
    .Y(_07002_)
  );
  sg13g2_o21ai_1 _16828_ (
    .A1(_02733_),
    .A2(_00021_),
    .B1(_03783_),
    .Y(_07003_)
  );
  sg13g2_a221oi_1 _16829_ (
    .A1(_00298_),
    .A2(_01191_),
    .B1(_07003_),
    .B2(_02287_),
    .C1(addr_i_8_),
    .Y(_07004_)
  );
  sg13g2_o21ai_1 _16830_ (
    .A1(addr_i_6_),
    .A2(_07002_),
    .B1(_07004_),
    .Y(_07006_)
  );
  sg13g2_a21oi_1 _16831_ (
    .A1(addr_i_2_),
    .A2(_02136_),
    .B1(_07790_),
    .Y(_07007_)
  );
  sg13g2_a22oi_1 _16832_ (
    .A1(_01160_),
    .A2(_01208_),
    .B1(_04778_),
    .B2(addr_i_6_),
    .Y(_07008_)
  );
  sg13g2_nor4_1 _16833_ (
    .A(_05888_),
    .B(_01194_),
    .C(_07007_),
    .D(_07008_),
    .Y(_07009_)
  );
  sg13g2_nor2_1 _16834_ (
    .A(_01658_),
    .B(_08951_),
    .Y(_07010_)
  );
  sg13g2_nor3_1 _16835_ (
    .A(addr_i_3_),
    .B(addr_i_4_),
    .C(_01054_),
    .Y(_07011_)
  );
  sg13g2_o21ai_1 _16836_ (
    .A1(_07010_),
    .A2(_07011_),
    .B1(addr_i_5_),
    .Y(_07012_)
  );
  sg13g2_nand3_1 _16837_ (
    .A(addr_i_7_),
    .B(_03669_),
    .C(_06571_),
    .Y(_07013_)
  );
  sg13g2_nand3_1 _16838_ (
    .A(_07009_),
    .B(_07012_),
    .C(_07013_),
    .Y(_07014_)
  );
  sg13g2_o21ai_1 _16839_ (
    .A1(_06999_),
    .A2(_07006_),
    .B1(_07014_),
    .Y(_07015_)
  );
  sg13g2_o21ai_1 _16840_ (
    .A1(addr_i_10_),
    .A2(_07015_),
    .B1(addr_i_9_),
    .Y(_07017_)
  );
  sg13g2_a21oi_1 _16841_ (
    .A1(addr_i_10_),
    .A2(_06996_),
    .B1(_07017_),
    .Y(_07018_)
  );
  sg13g2_nor2_1 _16842_ (
    .A(_09205_),
    .B(_00972_),
    .Y(_07019_)
  );
  sg13g2_o21ai_1 _16843_ (
    .A1(_02734_),
    .A2(_07019_),
    .B1(_03292_),
    .Y(_07020_)
  );
  sg13g2_o21ai_1 _16844_ (
    .A1(_03575_),
    .A2(_02578_),
    .B1(_07020_),
    .Y(_07021_)
  );
  sg13g2_a21oi_1 _16845_ (
    .A1(_00749_),
    .A2(_00531_),
    .B1(_07625_),
    .Y(_07022_)
  );
  sg13g2_a22oi_1 _16846_ (
    .A1(_01336_),
    .A2(_05542_),
    .B1(_07022_),
    .B2(_04837_),
    .Y(_07023_)
  );
  sg13g2_nor2_1 _16847_ (
    .A(_01391_),
    .B(_07023_),
    .Y(_07024_)
  );
  sg13g2_nor2_1 _16848_ (
    .A(addr_i_6_),
    .B(_00038_),
    .Y(_07025_)
  );
  sg13g2_nor2_1 _16849_ (
    .A(_07025_),
    .B(_01480_),
    .Y(_07026_)
  );
  sg13g2_a21oi_1 _16850_ (
    .A1(addr_i_6_),
    .A2(_04420_),
    .B1(addr_i_4_),
    .Y(_07028_)
  );
  sg13g2_a22oi_1 _16851_ (
    .A1(addr_i_4_),
    .A2(_07026_),
    .B1(_07028_),
    .B2(_03238_),
    .Y(_07029_)
  );
  sg13g2_a22oi_1 _16852_ (
    .A1(_00277_),
    .A2(_07021_),
    .B1(_07024_),
    .B2(_07029_),
    .Y(_07030_)
  );
  sg13g2_nand2_1 _16853_ (
    .A(_06740_),
    .B(_01302_),
    .Y(_07031_)
  );
  sg13g2_nand3_1 _16854_ (
    .A(addr_i_6_),
    .B(_00250_),
    .C(_07031_),
    .Y(_07032_)
  );
  sg13g2_a21oi_1 _16855_ (
    .A1(_00360_),
    .A2(_03854_),
    .B1(_00377_),
    .Y(_07033_)
  );
  sg13g2_nand2_1 _16856_ (
    .A(_02257_),
    .B(_07033_),
    .Y(_07034_)
  );
  sg13g2_a21oi_1 _16857_ (
    .A1(_00507_),
    .A2(_00105_),
    .B1(_00712_),
    .Y(_07035_)
  );
  sg13g2_a22oi_1 _16858_ (
    .A1(_07032_),
    .A2(_07034_),
    .B1(_03259_),
    .B2(_07035_),
    .Y(_07036_)
  );
  sg13g2_a21oi_1 _16859_ (
    .A1(_00476_),
    .A2(_01441_),
    .B1(_00116_),
    .Y(_07037_)
  );
  sg13g2_o21ai_1 _16860_ (
    .A1(_02215_),
    .A2(_07037_),
    .B1(addr_i_4_),
    .Y(_07039_)
  );
  sg13g2_nor4_1 _16861_ (
    .A(_01067_),
    .B(_01319_),
    .C(_00057_),
    .D(_05555_),
    .Y(_07040_)
  );
  sg13g2_nor3_1 _16862_ (
    .A(addr_i_3_),
    .B(_00644_),
    .C(_02069_),
    .Y(_07041_)
  );
  sg13g2_o21ai_1 _16863_ (
    .A1(_07040_),
    .A2(_07041_),
    .B1(_01008_),
    .Y(_07042_)
  );
  sg13g2_nand3_1 _16864_ (
    .A(addr_i_3_),
    .B(addr_i_7_),
    .C(_06132_),
    .Y(_07043_)
  );
  sg13g2_a21oi_1 _16865_ (
    .A1(_04451_),
    .A2(_07043_),
    .B1(_07337_),
    .Y(_07044_)
  );
  sg13g2_a21o_1 _16866_ (
    .A1(_06553_),
    .A2(_03943_),
    .B1(addr_i_5_),
    .X(_07045_)
  );
  sg13g2_a21oi_1 _16867_ (
    .A1(_03391_),
    .A2(_07045_),
    .B1(addr_i_7_),
    .Y(_07046_)
  );
  sg13g2_a22oi_1 _16868_ (
    .A1(addr_i_2_),
    .A2(_07042_),
    .B1(_07044_),
    .B2(_07046_),
    .Y(_07047_)
  );
  sg13g2_nor2_1 _16869_ (
    .A(addr_i_8_),
    .B(_07047_),
    .Y(_07048_)
  );
  sg13g2_a22oi_1 _16870_ (
    .A1(_07036_),
    .A2(_07039_),
    .B1(_07048_),
    .B2(_03841_),
    .Y(_07051_)
  );
  sg13g2_a22oi_1 _16871_ (
    .A1(_01774_),
    .A2(_07030_),
    .B1(_07051_),
    .B2(addr_i_9_),
    .Y(_07052_)
  );
  sg13g2_nor4_1 _16872_ (
    .A(addr_i_12_),
    .B(addr_i_11_),
    .C(_07018_),
    .D(_07052_),
    .Y(_07053_)
  );
  sg13g2_nor2_1 _16873_ (
    .A(_03540_),
    .B(_01197_),
    .Y(_07054_)
  );
  sg13g2_or2_1 _16874_ (
    .A(_02935_),
    .B(_07054_),
    .X(_07055_)
  );
  sg13g2_a21oi_1 _16875_ (
    .A1(addr_i_4_),
    .A2(_07055_),
    .B1(_01380_),
    .Y(_07056_)
  );
  sg13g2_o21ai_1 _16876_ (
    .A1(addr_i_6_),
    .A2(_07056_),
    .B1(_02577_),
    .Y(_07057_)
  );
  sg13g2_o21ai_1 _16877_ (
    .A1(_00087_),
    .A2(_06288_),
    .B1(addr_i_5_),
    .Y(_07058_)
  );
  sg13g2_o21ai_1 _16878_ (
    .A1(_00390_),
    .A2(_01216_),
    .B1(_07058_),
    .Y(_07059_)
  );
  sg13g2_a21oi_1 _16879_ (
    .A1(addr_i_4_),
    .A2(_04399_),
    .B1(_03150_),
    .Y(_07060_)
  );
  sg13g2_nor2_1 _16880_ (
    .A(_08266_),
    .B(_07060_),
    .Y(_07062_)
  );
  sg13g2_a221oi_1 _16881_ (
    .A1(_00169_),
    .A2(_01216_),
    .B1(_07059_),
    .B2(addr_i_3_),
    .C1(_07062_),
    .Y(_07063_)
  );
  sg13g2_a22oi_1 _16882_ (
    .A1(addr_i_2_),
    .A2(_01581_),
    .B1(_00242_),
    .B2(addr_i_3_),
    .Y(_07064_)
  );
  sg13g2_a22oi_1 _16883_ (
    .A1(_00591_),
    .A2(_02369_),
    .B1(_07064_),
    .B2(addr_i_4_),
    .Y(_07065_)
  );
  sg13g2_nand3_1 _16884_ (
    .A(addr_i_4_),
    .B(_00764_),
    .C(_02675_),
    .Y(_07066_)
  );
  sg13g2_nand2b_1 _16885_ (
    .A_N(_07065_),
    .B(_07066_),
    .Y(_07067_)
  );
  sg13g2_a22oi_1 _16886_ (
    .A1(_00239_),
    .A2(_09499_),
    .B1(_00645_),
    .B2(_01612_),
    .Y(_07068_)
  );
  sg13g2_nor2_1 _16887_ (
    .A(addr_i_3_),
    .B(_03466_),
    .Y(_07069_)
  );
  sg13g2_a22oi_1 _16888_ (
    .A1(addr_i_3_),
    .A2(_03467_),
    .B1(_07069_),
    .B2(_00396_),
    .Y(_07070_)
  );
  sg13g2_a21oi_1 _16889_ (
    .A1(_07067_),
    .A2(_07068_),
    .B1(_07070_),
    .Y(_07071_)
  );
  sg13g2_o21ai_1 _16890_ (
    .A1(_02368_),
    .A2(_07063_),
    .B1(_07071_),
    .Y(_07073_)
  );
  sg13g2_a221oi_1 _16891_ (
    .A1(_01350_),
    .A2(_07057_),
    .B1(_07073_),
    .B2(_01774_),
    .C1(_01359_),
    .Y(_07074_)
  );
  sg13g2_o21ai_1 _16892_ (
    .A1(_00597_),
    .A2(_01450_),
    .B1(_00386_),
    .Y(_07075_)
  );
  sg13g2_a21oi_1 _16893_ (
    .A1(addr_i_5_),
    .A2(_01103_),
    .B1(_02136_),
    .Y(_07076_)
  );
  sg13g2_o21ai_1 _16894_ (
    .A1(_00474_),
    .A2(_07076_),
    .B1(addr_i_2_),
    .Y(_07077_)
  );
  sg13g2_nand3_1 _16895_ (
    .A(_00782_),
    .B(_07075_),
    .C(_07077_),
    .Y(_07078_)
  );
  sg13g2_a21oi_1 _16896_ (
    .A1(_09260_),
    .A2(_00405_),
    .B1(addr_i_3_),
    .Y(_07079_)
  );
  sg13g2_a21oi_1 _16897_ (
    .A1(_01257_),
    .A2(_00434_),
    .B1(_01144_),
    .Y(_07080_)
  );
  sg13g2_a22oi_1 _16898_ (
    .A1(_01191_),
    .A2(_01555_),
    .B1(_07079_),
    .B2(_07080_),
    .Y(_07081_)
  );
  sg13g2_nor2_1 _16899_ (
    .A(_01630_),
    .B(_07081_),
    .Y(_07082_)
  );
  sg13g2_nor3_1 _16900_ (
    .A(addr_i_5_),
    .B(_09492_),
    .C(_02268_),
    .Y(_07084_)
  );
  sg13g2_a21oi_1 _16901_ (
    .A1(_00377_),
    .A2(_00409_),
    .B1(_07084_),
    .Y(_07085_)
  );
  sg13g2_o21ai_1 _16902_ (
    .A1(_00377_),
    .A2(_03150_),
    .B1(_02344_),
    .Y(_07086_)
  );
  sg13g2_nand2_1 _16903_ (
    .A(addr_i_3_),
    .B(_01252_),
    .Y(_07087_)
  );
  sg13g2_a21oi_1 _16904_ (
    .A1(_02063_),
    .A2(_02437_),
    .B1(_07087_),
    .Y(_07088_)
  );
  sg13g2_a21oi_1 _16905_ (
    .A1(_01290_),
    .A2(_00434_),
    .B1(addr_i_4_),
    .Y(_07089_)
  );
  sg13g2_o21ai_1 _16906_ (
    .A1(_00080_),
    .A2(_01222_),
    .B1(addr_i_8_),
    .Y(_07090_)
  );
  sg13g2_a22oi_1 _16907_ (
    .A1(_07086_),
    .A2(_07088_),
    .B1(_07089_),
    .B2(_07090_),
    .Y(_07091_)
  );
  sg13g2_o21ai_1 _16908_ (
    .A1(addr_i_3_),
    .A2(_07085_),
    .B1(_07091_),
    .Y(_07092_)
  );
  sg13g2_o21ai_1 _16909_ (
    .A1(_07078_),
    .A2(_07082_),
    .B1(_07092_),
    .Y(_07093_)
  );
  sg13g2_a21oi_1 _16910_ (
    .A1(addr_i_6_),
    .A2(_02472_),
    .B1(addr_i_3_),
    .Y(_07095_)
  );
  sg13g2_o21ai_1 _16911_ (
    .A1(_01500_),
    .A2(_07095_),
    .B1(addr_i_5_),
    .Y(_07096_)
  );
  sg13g2_o21ai_1 _16912_ (
    .A1(_00305_),
    .A2(_02542_),
    .B1(addr_i_3_),
    .Y(_07097_)
  );
  sg13g2_nand3_1 _16913_ (
    .A(_05780_),
    .B(_07096_),
    .C(_07097_),
    .Y(_07098_)
  );
  sg13g2_nor2_1 _16914_ (
    .A(_08431_),
    .B(_07558_),
    .Y(_07099_)
  );
  sg13g2_o21ai_1 _16915_ (
    .A1(_00598_),
    .A2(_07099_),
    .B1(addr_i_4_),
    .Y(_07100_)
  );
  sg13g2_a21oi_1 _16916_ (
    .A1(_01168_),
    .A2(_07100_),
    .B1(_03238_),
    .Y(_07101_)
  );
  sg13g2_a21oi_1 _16917_ (
    .A1(_01119_),
    .A2(_07098_),
    .B1(_07101_),
    .Y(_07102_)
  );
  sg13g2_nand2_1 _16918_ (
    .A(_00403_),
    .B(_03267_),
    .Y(_07103_)
  );
  sg13g2_o21ai_1 _16919_ (
    .A1(_02513_),
    .A2(_03077_),
    .B1(_07103_),
    .Y(_07104_)
  );
  sg13g2_o21ai_1 _16920_ (
    .A1(_00401_),
    .A2(_02486_),
    .B1(addr_i_6_),
    .Y(_07106_)
  );
  sg13g2_a21oi_1 _16921_ (
    .A1(_03871_),
    .A2(_07106_),
    .B1(_03062_),
    .Y(_07107_)
  );
  sg13g2_a22oi_1 _16922_ (
    .A1(_00440_),
    .A2(_07104_),
    .B1(_07107_),
    .B2(addr_i_9_),
    .Y(_07108_)
  );
  sg13g2_a221oi_1 _16923_ (
    .A1(addr_i_9_),
    .A2(_07093_),
    .B1(_07102_),
    .B2(_07108_),
    .C1(addr_i_10_),
    .Y(_07109_)
  );
  sg13g2_a21o_1 _16924_ (
    .A1(_04442_),
    .A2(_01179_),
    .B1(_00012_),
    .X(_07110_)
  );
  sg13g2_nand3_1 _16925_ (
    .A(_01892_),
    .B(_01268_),
    .C(_04745_),
    .Y(_07111_)
  );
  sg13g2_nand3_1 _16926_ (
    .A(addr_i_7_),
    .B(_00150_),
    .C(_09479_),
    .Y(_07112_)
  );
  sg13g2_nand3_1 _16927_ (
    .A(_05218_),
    .B(_01872_),
    .C(_01795_),
    .Y(_07113_)
  );
  sg13g2_nand3_1 _16928_ (
    .A(addr_i_4_),
    .B(_07112_),
    .C(_07113_),
    .Y(_07114_)
  );
  sg13g2_o21ai_1 _16929_ (
    .A1(_00400_),
    .A2(_02376_),
    .B1(addr_i_7_),
    .Y(_07115_)
  );
  sg13g2_nor2_1 _16930_ (
    .A(_05711_),
    .B(_02638_),
    .Y(_07117_)
  );
  sg13g2_nor2_1 _16931_ (
    .A(_06950_),
    .B(_07117_),
    .Y(_07118_)
  );
  sg13g2_mux2_1 _16932_ (
    .A0(_07115_),
    .A1(_07118_),
    .S(_02287_),
    .X(_07119_)
  );
  sg13g2_nand3_1 _16933_ (
    .A(addr_i_6_),
    .B(_07114_),
    .C(_07119_),
    .Y(_07120_)
  );
  sg13g2_nand4_1 _16934_ (
    .A(addr_i_8_),
    .B(_07110_),
    .C(_07111_),
    .D(_07120_),
    .Y(_07121_)
  );
  sg13g2_nand3_1 _16935_ (
    .A(addr_i_2_),
    .B(_00151_),
    .C(_01060_),
    .Y(_07122_)
  );
  sg13g2_nand3_1 _16936_ (
    .A(_08011_),
    .B(_03226_),
    .C(_03669_),
    .Y(_07123_)
  );
  sg13g2_nor2_1 _16937_ (
    .A(_05921_),
    .B(_01144_),
    .Y(_07124_)
  );
  sg13g2_a21oi_1 _16938_ (
    .A1(_07122_),
    .A2(_07123_),
    .B1(_07124_),
    .Y(_07125_)
  );
  sg13g2_nand3_1 _16939_ (
    .A(_00228_),
    .B(_09478_),
    .C(_06909_),
    .Y(_07126_)
  );
  sg13g2_a21oi_1 _16940_ (
    .A1(_00762_),
    .A2(_02002_),
    .B1(_00507_),
    .Y(_07128_)
  );
  sg13g2_a22oi_1 _16941_ (
    .A1(_00169_),
    .A2(_07126_),
    .B1(_07128_),
    .B2(addr_i_8_),
    .Y(_07129_)
  );
  sg13g2_o21ai_1 _16942_ (
    .A1(addr_i_7_),
    .A2(_07125_),
    .B1(_07129_),
    .Y(_07130_)
  );
  sg13g2_and3_1 _16943_ (
    .A(_01176_),
    .B(_07121_),
    .C(_07130_),
    .X(_07131_)
  );
  sg13g2_o21ai_1 _16944_ (
    .A1(_01227_),
    .A2(_02161_),
    .B1(addr_i_2_),
    .Y(_07132_)
  );
  sg13g2_o21ai_1 _16945_ (
    .A1(_01616_),
    .A2(_01480_),
    .B1(_00123_),
    .Y(_07133_)
  );
  sg13g2_nand3_1 _16946_ (
    .A(_00403_),
    .B(_07132_),
    .C(_07133_),
    .Y(_07134_)
  );
  sg13g2_nor3_1 _16947_ (
    .A(_07889_),
    .B(_08575_),
    .C(_03360_),
    .Y(_07135_)
  );
  sg13g2_nand4_1 _16948_ (
    .A(_01892_),
    .B(_00651_),
    .C(_08022_),
    .D(_06067_),
    .Y(_07136_)
  );
  sg13g2_o21ai_1 _16949_ (
    .A1(_00053_),
    .A2(_07135_),
    .B1(_07136_),
    .Y(_07137_)
  );
  sg13g2_a22oi_1 _16950_ (
    .A1(_05834_),
    .A2(_07134_),
    .B1(_07137_),
    .B2(_00114_),
    .Y(_07139_)
  );
  sg13g2_nand2_1 _16951_ (
    .A(_03431_),
    .B(_01872_),
    .Y(_07140_)
  );
  sg13g2_a22oi_1 _16952_ (
    .A1(_01794_),
    .A2(_07140_),
    .B1(_03164_),
    .B2(_00227_),
    .Y(_07141_)
  );
  sg13g2_nor2_1 _16953_ (
    .A(_00390_),
    .B(_07141_),
    .Y(_07142_)
  );
  sg13g2_nand3_1 _16954_ (
    .A(_07337_),
    .B(_09487_),
    .C(_02028_),
    .Y(_07143_)
  );
  sg13g2_a21oi_1 _16955_ (
    .A1(_00827_),
    .A2(_01355_),
    .B1(_07143_),
    .Y(_07144_)
  );
  sg13g2_o21ai_1 _16956_ (
    .A1(addr_i_2_),
    .A2(_02342_),
    .B1(_02467_),
    .Y(_07145_)
  );
  sg13g2_a21oi_1 _16957_ (
    .A1(_00371_),
    .A2(_05012_),
    .B1(_00191_),
    .Y(_07146_)
  );
  sg13g2_a22oi_1 _16958_ (
    .A1(_00048_),
    .A2(_07145_),
    .B1(_07146_),
    .B2(_04767_),
    .Y(_07147_)
  );
  sg13g2_nor4_1 _16959_ (
    .A(addr_i_8_),
    .B(_07142_),
    .C(_07144_),
    .D(_07147_),
    .Y(_07148_)
  );
  sg13g2_nor3_1 _16960_ (
    .A(_00109_),
    .B(_07139_),
    .C(_07148_),
    .Y(_07150_)
  );
  sg13g2_nor4_1 _16961_ (
    .A(_01451_),
    .B(_07109_),
    .C(_07131_),
    .D(_07150_),
    .Y(_07151_)
  );
  sg13g2_nor4_1 _16962_ (
    .A(_06979_),
    .B(_07053_),
    .C(_07074_),
    .D(_07151_),
    .Y(data_o_2_)
  );
  sg13g2_o21ai_1 _16963_ (
    .A1(addr_i_5_),
    .A2(_04371_),
    .B1(_02694_),
    .Y(_07152_)
  );
  sg13g2_nand3_1 _16964_ (
    .A(addr_i_3_),
    .B(_01983_),
    .C(_02032_),
    .Y(_07153_)
  );
  sg13g2_o21ai_1 _16965_ (
    .A1(addr_i_3_),
    .A2(_07152_),
    .B1(_07153_),
    .Y(_07154_)
  );
  sg13g2_nand3_1 _16966_ (
    .A(_02165_),
    .B(_01518_),
    .C(_07154_),
    .Y(_07155_)
  );
  sg13g2_a21oi_1 _16967_ (
    .A1(addr_i_3_),
    .A2(_01085_),
    .B1(_09172_),
    .Y(_07156_)
  );
  sg13g2_nand2_1 _16968_ (
    .A(_09393_),
    .B(_08254_),
    .Y(_07157_)
  );
  sg13g2_a21oi_1 _16969_ (
    .A1(addr_i_4_),
    .A2(_07157_),
    .B1(_01622_),
    .Y(_07158_)
  );
  sg13g2_a21oi_1 _16970_ (
    .A1(_00117_),
    .A2(_05430_),
    .B1(_05379_),
    .Y(_07161_)
  );
  sg13g2_a21oi_1 _16971_ (
    .A1(_06077_),
    .A2(_01960_),
    .B1(_03270_),
    .Y(_07162_)
  );
  sg13g2_nor2_1 _16972_ (
    .A(addr_i_4_),
    .B(_07162_),
    .Y(_07163_)
  );
  sg13g2_a22oi_1 _16973_ (
    .A1(addr_i_4_),
    .A2(_07161_),
    .B1(_07163_),
    .B2(addr_i_7_),
    .Y(_07164_)
  );
  sg13g2_a21oi_1 _16974_ (
    .A1(_07156_),
    .A2(_07158_),
    .B1(_07164_),
    .Y(_07165_)
  );
  sg13g2_a22oi_1 _16975_ (
    .A1(_00210_),
    .A2(_00514_),
    .B1(_03137_),
    .B2(_03267_),
    .Y(_07166_)
  );
  sg13g2_nand3b_1 _16976_ (
    .A_N(_00839_),
    .B(_06779_),
    .C(_07166_),
    .Y(_07167_)
  );
  sg13g2_nand2_1 _16977_ (
    .A(_02141_),
    .B(_00828_),
    .Y(_07168_)
  );
  sg13g2_a21oi_1 _16978_ (
    .A1(_06508_),
    .A2(_07168_),
    .B1(_02213_),
    .Y(_07169_)
  );
  sg13g2_a21oi_1 _16979_ (
    .A1(_00872_),
    .A2(_01245_),
    .B1(_02294_),
    .Y(_07170_)
  );
  sg13g2_a22oi_1 _16980_ (
    .A1(addr_i_7_),
    .A2(_07167_),
    .B1(_07169_),
    .B2(_07170_),
    .Y(_07172_)
  );
  sg13g2_nor2_1 _16981_ (
    .A(_00014_),
    .B(_02055_),
    .Y(_07173_)
  );
  sg13g2_a21oi_1 _16982_ (
    .A1(_04318_),
    .A2(_03139_),
    .B1(_04265_),
    .Y(_07174_)
  );
  sg13g2_o21ai_1 _16983_ (
    .A1(addr_i_3_),
    .A2(_07173_),
    .B1(_07174_),
    .Y(_07175_)
  );
  sg13g2_o21ai_1 _16984_ (
    .A1(_03523_),
    .A2(_07175_),
    .B1(_05218_),
    .Y(_07176_)
  );
  sg13g2_nor2_1 _16985_ (
    .A(_00824_),
    .B(_01782_),
    .Y(_07177_)
  );
  sg13g2_a22oi_1 _16986_ (
    .A1(_00199_),
    .A2(_01552_),
    .B1(_01582_),
    .B2(_00839_),
    .Y(_07178_)
  );
  sg13g2_nand4_1 _16987_ (
    .A(_03205_),
    .B(_01168_),
    .C(_07177_),
    .D(_07178_),
    .Y(_07179_)
  );
  sg13g2_a21oi_1 _16988_ (
    .A1(_01252_),
    .A2(_02920_),
    .B1(_00719_),
    .Y(_07180_)
  );
  sg13g2_a221oi_1 _16989_ (
    .A1(_01202_),
    .A2(_09498_),
    .B1(_07179_),
    .B2(addr_i_7_),
    .C1(_07180_),
    .Y(_07181_)
  );
  sg13g2_mux4_1 _16990_ (
    .A0(_07165_),
    .A1(_07172_),
    .A2(_07176_),
    .A3(_07181_),
    .S0(addr_i_8_),
    .S1(_09315_),
    .X(_07183_)
  );
  sg13g2_nand2_1 _16991_ (
    .A(_07155_),
    .B(_07183_),
    .Y(_07184_)
  );
  sg13g2_o21ai_1 _16992_ (
    .A1(_06607_),
    .A2(_00635_),
    .B1(_00293_),
    .Y(_07185_)
  );
  sg13g2_o21ai_1 _16993_ (
    .A1(_00115_),
    .A2(_01437_),
    .B1(_07185_),
    .Y(_07186_)
  );
  sg13g2_nor2_1 _16994_ (
    .A(addr_i_4_),
    .B(_01147_),
    .Y(_07187_)
  );
  sg13g2_a22oi_1 _16995_ (
    .A1(addr_i_4_),
    .A2(_07186_),
    .B1(_07187_),
    .B2(_02652_),
    .Y(_07188_)
  );
  sg13g2_nand2_1 _16996_ (
    .A(_02427_),
    .B(_05255_),
    .Y(_07189_)
  );
  sg13g2_o21ai_1 _16997_ (
    .A1(_05280_),
    .A2(_09498_),
    .B1(addr_i_2_),
    .Y(_07190_)
  );
  sg13g2_o21ai_1 _16998_ (
    .A1(addr_i_5_),
    .A2(_00294_),
    .B1(_02462_),
    .Y(_07191_)
  );
  sg13g2_a21oi_1 _16999_ (
    .A1(_07190_),
    .A2(_07191_),
    .B1(addr_i_4_),
    .Y(_07192_)
  );
  sg13g2_a22oi_1 _17000_ (
    .A1(addr_i_4_),
    .A2(_07189_),
    .B1(_07192_),
    .B2(_00113_),
    .Y(_07194_)
  );
  sg13g2_o21ai_1 _17001_ (
    .A1(addr_i_2_),
    .A2(_07188_),
    .B1(_07194_),
    .Y(_07195_)
  );
  sg13g2_o21ai_1 _17002_ (
    .A1(addr_i_4_),
    .A2(_01413_),
    .B1(_01070_),
    .Y(_07196_)
  );
  sg13g2_o21ai_1 _17003_ (
    .A1(_00001_),
    .A2(_00294_),
    .B1(addr_i_3_),
    .Y(_07197_)
  );
  sg13g2_a21oi_1 _17004_ (
    .A1(_00994_),
    .A2(_07197_),
    .B1(addr_i_6_),
    .Y(_07198_)
  );
  sg13g2_o21ai_1 _17005_ (
    .A1(_00534_),
    .A2(_03648_),
    .B1(addr_i_7_),
    .Y(_07199_)
  );
  sg13g2_nand2_1 _17006_ (
    .A(_07282_),
    .B(_07199_),
    .Y(_07200_)
  );
  sg13g2_a22oi_1 _17007_ (
    .A1(_00223_),
    .A2(_07196_),
    .B1(_07198_),
    .B2(_07200_),
    .Y(_07201_)
  );
  sg13g2_a21oi_1 _17008_ (
    .A1(_02529_),
    .A2(_01463_),
    .B1(addr_i_7_),
    .Y(_07202_)
  );
  sg13g2_a21oi_1 _17009_ (
    .A1(_00358_),
    .A2(_01234_),
    .B1(_00083_),
    .Y(_07203_)
  );
  sg13g2_o21ai_1 _17010_ (
    .A1(_07202_),
    .A2(_07203_),
    .B1(addr_i_5_),
    .Y(_07205_)
  );
  sg13g2_a21oi_1 _17011_ (
    .A1(_07201_),
    .A2(_07205_),
    .B1(_04705_),
    .Y(_07206_)
  );
  sg13g2_a21oi_1 _17012_ (
    .A1(_00284_),
    .A2(_08221_),
    .B1(_00498_),
    .Y(_07207_)
  );
  sg13g2_a21oi_1 _17013_ (
    .A1(_01077_),
    .A2(_03167_),
    .B1(_00961_),
    .Y(_07208_)
  );
  sg13g2_o21ai_1 _17014_ (
    .A1(_07207_),
    .A2(_07208_),
    .B1(addr_i_5_),
    .Y(_07209_)
  );
  sg13g2_o21ai_1 _17015_ (
    .A1(addr_i_2_),
    .A2(_06927_),
    .B1(_00474_),
    .Y(_07210_)
  );
  sg13g2_o21ai_1 _17016_ (
    .A1(_02698_),
    .A2(_03562_),
    .B1(_05218_),
    .Y(_07211_)
  );
  sg13g2_nor3_1 _17017_ (
    .A(_05070_),
    .B(_06398_),
    .C(_02470_),
    .Y(_07212_)
  );
  sg13g2_o21ai_1 _17018_ (
    .A1(_01093_),
    .A2(_07212_),
    .B1(_00083_),
    .Y(_07213_)
  );
  sg13g2_nand4_1 _17019_ (
    .A(_07209_),
    .B(_07210_),
    .C(_07211_),
    .D(_07213_),
    .Y(_07214_)
  );
  sg13g2_a22oi_1 _17020_ (
    .A1(_02467_),
    .A2(_02690_),
    .B1(_01279_),
    .B2(_00802_),
    .Y(_07216_)
  );
  sg13g2_a221oi_1 _17021_ (
    .A1(_00960_),
    .A2(_09348_),
    .B1(_07168_),
    .B2(addr_i_6_),
    .C1(_07603_),
    .Y(_07217_)
  );
  sg13g2_or2_1 _17022_ (
    .A(addr_i_9_),
    .B(_07217_),
    .X(_07218_)
  );
  sg13g2_a22oi_1 _17023_ (
    .A1(addr_i_8_),
    .A2(_07214_),
    .B1(_07216_),
    .B2(_07218_),
    .Y(_07219_)
  );
  sg13g2_a22oi_1 _17024_ (
    .A1(_07195_),
    .A2(_07206_),
    .B1(_07219_),
    .B2(addr_i_10_),
    .Y(_07220_)
  );
  sg13g2_a22oi_1 _17025_ (
    .A1(addr_i_10_),
    .A2(_07184_),
    .B1(_07220_),
    .B2(addr_i_11_),
    .Y(_07221_)
  );
  sg13g2_nand2_1 _17026_ (
    .A(_08564_),
    .B(_03314_),
    .Y(_07222_)
  );
  sg13g2_nor2_1 _17027_ (
    .A(_00927_),
    .B(_07222_),
    .Y(_07223_)
  );
  sg13g2_a221oi_1 _17028_ (
    .A1(addr_i_5_),
    .A2(_02200_),
    .B1(_02785_),
    .B2(addr_i_7_),
    .C1(_07223_),
    .Y(_07224_)
  );
  sg13g2_a21oi_1 _17029_ (
    .A1(_08376_),
    .A2(_00965_),
    .B1(_06176_),
    .Y(_07225_)
  );
  sg13g2_a21oi_1 _17030_ (
    .A1(_08410_),
    .A2(_02638_),
    .B1(_07225_),
    .Y(_07227_)
  );
  sg13g2_a21oi_1 _17031_ (
    .A1(_09509_),
    .A2(_00158_),
    .B1(_02990_),
    .Y(_07228_)
  );
  sg13g2_nand2_1 _17032_ (
    .A(_07227_),
    .B(_07228_),
    .Y(_07229_)
  );
  sg13g2_o21ai_1 _17033_ (
    .A1(addr_i_3_),
    .A2(_07224_),
    .B1(_07229_),
    .Y(_07230_)
  );
  sg13g2_a21oi_1 _17034_ (
    .A1(_01301_),
    .A2(_02529_),
    .B1(addr_i_3_),
    .Y(_07231_)
  );
  sg13g2_o21ai_1 _17035_ (
    .A1(_08343_),
    .A2(_01086_),
    .B1(addr_i_3_),
    .Y(_07232_)
  );
  sg13g2_nand3_1 _17036_ (
    .A(addr_i_7_),
    .B(_05780_),
    .C(_07232_),
    .Y(_07233_)
  );
  sg13g2_a21oi_1 _17037_ (
    .A1(_03665_),
    .A2(_00890_),
    .B1(_03106_),
    .Y(_07234_)
  );
  sg13g2_o21ai_1 _17038_ (
    .A1(addr_i_6_),
    .A2(_01472_),
    .B1(_00635_),
    .Y(_07235_)
  );
  sg13g2_o21ai_1 _17039_ (
    .A1(addr_i_7_),
    .A2(_07234_),
    .B1(_07235_),
    .Y(_07236_)
  );
  sg13g2_a21oi_1 _17040_ (
    .A1(_03875_),
    .A2(_02319_),
    .B1(_00441_),
    .Y(_07238_)
  );
  sg13g2_a22oi_1 _17041_ (
    .A1(addr_i_5_),
    .A2(_07236_),
    .B1(_07238_),
    .B2(_05888_),
    .Y(_07239_)
  );
  sg13g2_o21ai_1 _17042_ (
    .A1(_07231_),
    .A2(_07233_),
    .B1(_07239_),
    .Y(_07240_)
  );
  sg13g2_o21ai_1 _17043_ (
    .A1(addr_i_8_),
    .A2(_07230_),
    .B1(_07240_),
    .Y(_07241_)
  );
  sg13g2_a221oi_1 _17044_ (
    .A1(_00294_),
    .A2(_02383_),
    .B1(_00578_),
    .B2(addr_i_5_),
    .C1(_01867_),
    .Y(_07242_)
  );
  sg13g2_o21ai_1 _17045_ (
    .A1(_01113_),
    .A2(_00098_),
    .B1(_00878_),
    .Y(_07243_)
  );
  sg13g2_nand2_1 _17046_ (
    .A(_00445_),
    .B(_07243_),
    .Y(_07244_)
  );
  sg13g2_a21o_1 _17047_ (
    .A1(_07242_),
    .A2(_07244_),
    .B1(addr_i_3_),
    .X(_07245_)
  );
  sg13g2_o21ai_1 _17048_ (
    .A1(_04196_),
    .A2(_04915_),
    .B1(_04108_),
    .Y(_07246_)
  );
  sg13g2_o21ai_1 _17049_ (
    .A1(_09509_),
    .A2(_05757_),
    .B1(_07246_),
    .Y(_07247_)
  );
  sg13g2_nor3_1 _17050_ (
    .A(_01065_),
    .B(_01024_),
    .C(_01015_),
    .Y(_07249_)
  );
  sg13g2_a22oi_1 _17051_ (
    .A1(addr_i_3_),
    .A2(_07247_),
    .B1(_07249_),
    .B2(addr_i_8_),
    .Y(_07250_)
  );
  sg13g2_o21ai_1 _17052_ (
    .A1(addr_i_3_),
    .A2(_02173_),
    .B1(_00024_),
    .Y(_07251_)
  );
  sg13g2_a21oi_1 _17053_ (
    .A1(_03743_),
    .A2(_01182_),
    .B1(_08332_),
    .Y(_07252_)
  );
  sg13g2_a22oi_1 _17054_ (
    .A1(addr_i_3_),
    .A2(_06643_),
    .B1(_07251_),
    .B2(_07252_),
    .Y(_07253_)
  );
  sg13g2_a22oi_1 _17055_ (
    .A1(_00050_),
    .A2(_01337_),
    .B1(addr_i_3_),
    .B2(_05302_),
    .Y(_07254_)
  );
  sg13g2_a21oi_1 _17056_ (
    .A1(_09149_),
    .A2(_02089_),
    .B1(_00549_),
    .Y(_07255_)
  );
  sg13g2_a22oi_1 _17057_ (
    .A1(_00594_),
    .A2(_09499_),
    .B1(_07254_),
    .B2(_07255_),
    .Y(_07256_)
  );
  sg13g2_o21ai_1 _17058_ (
    .A1(addr_i_4_),
    .A2(_07253_),
    .B1(_07256_),
    .Y(_07257_)
  );
  sg13g2_a221oi_1 _17059_ (
    .A1(_07245_),
    .A2(_07250_),
    .B1(_07257_),
    .B2(addr_i_8_),
    .C1(addr_i_9_),
    .Y(_07258_)
  );
  sg13g2_a22oi_1 _17060_ (
    .A1(addr_i_9_),
    .A2(_07241_),
    .B1(_07258_),
    .B2(addr_i_10_),
    .Y(_07260_)
  );
  sg13g2_mux2_1 _17061_ (
    .A0(_00786_),
    .A1(_04613_),
    .S(_00593_),
    .X(_07261_)
  );
  sg13g2_o21ai_1 _17062_ (
    .A1(_01402_),
    .A2(_07261_),
    .B1(addr_i_2_),
    .Y(_07262_)
  );
  sg13g2_a21o_1 _17063_ (
    .A1(_04662_),
    .A2(_04252_),
    .B1(_00692_),
    .X(_07263_)
  );
  sg13g2_a21oi_1 _17064_ (
    .A1(_07262_),
    .A2(_07263_),
    .B1(_01099_),
    .Y(_07264_)
  );
  sg13g2_nand2_1 _17065_ (
    .A(_01257_),
    .B(_00595_),
    .Y(_07265_)
  );
  sg13g2_o21ai_1 _17066_ (
    .A1(addr_i_5_),
    .A2(_00304_),
    .B1(addr_i_2_),
    .Y(_07266_)
  );
  sg13g2_a21oi_1 _17067_ (
    .A1(_01224_),
    .A2(_07266_),
    .B1(_05867_),
    .Y(_07267_)
  );
  sg13g2_a22oi_1 _17068_ (
    .A1(addr_i_4_),
    .A2(_07265_),
    .B1(_07267_),
    .B2(_00588_),
    .Y(_07268_)
  );
  sg13g2_nand2_1 _17069_ (
    .A(_01370_),
    .B(_03108_),
    .Y(_07269_)
  );
  sg13g2_a22oi_1 _17070_ (
    .A1(addr_i_3_),
    .A2(_07269_),
    .B1(_01582_),
    .B2(_09359_),
    .Y(_07272_)
  );
  sg13g2_o21ai_1 _17071_ (
    .A1(_00484_),
    .A2(_03401_),
    .B1(_01051_),
    .Y(_07273_)
  );
  sg13g2_o21ai_1 _17072_ (
    .A1(_02634_),
    .A2(_02289_),
    .B1(_00429_),
    .Y(_07274_)
  );
  sg13g2_a21o_1 _17073_ (
    .A1(addr_i_3_),
    .A2(_07273_),
    .B1(_07274_),
    .X(_07275_)
  );
  sg13g2_o21ai_1 _17074_ (
    .A1(_01285_),
    .A2(_07272_),
    .B1(_07275_),
    .Y(_07276_)
  );
  sg13g2_nor4_1 _17075_ (
    .A(addr_i_9_),
    .B(_07264_),
    .C(_07268_),
    .D(_07276_),
    .Y(_07277_)
  );
  sg13g2_a22oi_1 _17076_ (
    .A1(addr_i_2_),
    .A2(_03336_),
    .B1(_02441_),
    .B2(addr_i_3_),
    .Y(_07278_)
  );
  sg13g2_nand3_1 _17077_ (
    .A(addr_i_3_),
    .B(_00371_),
    .C(_00228_),
    .Y(_07279_)
  );
  sg13g2_nand3b_1 _17078_ (
    .A_N(_07278_),
    .B(_07279_),
    .C(addr_i_7_),
    .Y(_07280_)
  );
  sg13g2_o21ai_1 _17079_ (
    .A1(_01033_),
    .A2(_00950_),
    .B1(_06132_),
    .Y(_07281_)
  );
  sg13g2_a21oi_1 _17080_ (
    .A1(_05745_),
    .A2(_08464_),
    .B1(_00927_),
    .Y(_07283_)
  );
  sg13g2_nand2_1 _17081_ (
    .A(_02053_),
    .B(_07812_),
    .Y(_07284_)
  );
  sg13g2_a21oi_1 _17082_ (
    .A1(addr_i_5_),
    .A2(_07284_),
    .B1(_03167_),
    .Y(_07285_)
  );
  sg13g2_a22oi_1 _17083_ (
    .A1(_01308_),
    .A2(_07281_),
    .B1(_07283_),
    .B2(_07285_),
    .Y(_07286_)
  );
  sg13g2_a21oi_1 _17084_ (
    .A1(_07280_),
    .A2(_07286_),
    .B1(addr_i_8_),
    .Y(_07287_)
  );
  sg13g2_nand2_1 _17085_ (
    .A(_05966_),
    .B(_02645_),
    .Y(_07288_)
  );
  sg13g2_nand2_1 _17086_ (
    .A(_03106_),
    .B(_01197_),
    .Y(_07289_)
  );
  sg13g2_nand3_1 _17087_ (
    .A(addr_i_2_),
    .B(_07288_),
    .C(_07289_),
    .Y(_07290_)
  );
  sg13g2_nand3_1 _17088_ (
    .A(_00593_),
    .B(_04362_),
    .C(_02020_),
    .Y(_07291_)
  );
  sg13g2_nand3_1 _17089_ (
    .A(_02343_),
    .B(_04765_),
    .C(_07291_),
    .Y(_07292_)
  );
  sg13g2_a21o_1 _17090_ (
    .A1(_07290_),
    .A2(_07292_),
    .B1(_01011_),
    .X(_07294_)
  );
  sg13g2_o21ai_1 _17091_ (
    .A1(_00557_),
    .A2(_01375_),
    .B1(_02387_),
    .Y(_07295_)
  );
  sg13g2_o21ai_1 _17092_ (
    .A1(_06298_),
    .A2(_01436_),
    .B1(addr_i_3_),
    .Y(_07296_)
  );
  sg13g2_nand4_1 _17093_ (
    .A(_01589_),
    .B(_07934_),
    .C(_07295_),
    .D(_07296_),
    .Y(_07297_)
  );
  sg13g2_nand3_1 _17094_ (
    .A(addr_i_9_),
    .B(_07294_),
    .C(_07297_),
    .Y(_07298_)
  );
  sg13g2_o21ai_1 _17095_ (
    .A1(_07287_),
    .A2(_07298_),
    .B1(addr_i_10_),
    .Y(_07299_)
  );
  sg13g2_o21ai_1 _17096_ (
    .A1(_07277_),
    .A2(_07299_),
    .B1(addr_i_11_),
    .Y(_07300_)
  );
  sg13g2_o21ai_1 _17097_ (
    .A1(_07260_),
    .A2(_07300_),
    .B1(_02996_),
    .Y(_07301_)
  );
  sg13g2_nor2_1 _17098_ (
    .A(_07221_),
    .B(_07301_),
    .Y(_07302_)
  );
  sg13g2_nor2_1 _17099_ (
    .A(_00827_),
    .B(_03993_),
    .Y(_07303_)
  );
  sg13g2_o21ai_1 _17100_ (
    .A1(addr_i_4_),
    .A2(_07303_),
    .B1(_05490_),
    .Y(_07305_)
  );
  sg13g2_o21ai_1 _17101_ (
    .A1(_02578_),
    .A2(_08232_),
    .B1(_00113_),
    .Y(_07306_)
  );
  sg13g2_nand3_1 _17102_ (
    .A(_05247_),
    .B(_00884_),
    .C(_03324_),
    .Y(_07307_)
  );
  sg13g2_a21oi_1 _17103_ (
    .A1(_00056_),
    .A2(_07307_),
    .B1(addr_i_2_),
    .Y(_07308_)
  );
  sg13g2_a22oi_1 _17104_ (
    .A1(_09474_),
    .A2(_07305_),
    .B1(_07306_),
    .B2(_07308_),
    .Y(_07309_)
  );
  sg13g2_o21ai_1 _17105_ (
    .A1(_08144_),
    .A2(_02424_),
    .B1(_05711_),
    .Y(_07310_)
  );
  sg13g2_nand2_1 _17106_ (
    .A(_05819_),
    .B(_07310_),
    .Y(_07311_)
  );
  sg13g2_a21oi_1 _17107_ (
    .A1(_02930_),
    .A2(_04200_),
    .B1(addr_i_3_),
    .Y(_07312_)
  );
  sg13g2_a21oi_1 _17108_ (
    .A1(addr_i_6_),
    .A2(_07311_),
    .B1(_07312_),
    .Y(_07313_)
  );
  sg13g2_o21ai_1 _17109_ (
    .A1(addr_i_7_),
    .A2(_07313_),
    .B1(_03448_),
    .Y(_07314_)
  );
  sg13g2_nor2b_1 _17110_ (
    .A(_07309_),
    .B_N(_07314_),
    .Y(_07316_)
  );
  sg13g2_o21ai_1 _17111_ (
    .A1(addr_i_9_),
    .A2(_07316_),
    .B1(_02036_),
    .Y(_07317_)
  );
  sg13g2_nor2_1 _17112_ (
    .A(_01240_),
    .B(_00807_),
    .Y(_07318_)
  );
  sg13g2_o21ai_1 _17113_ (
    .A1(_01634_),
    .A2(_02033_),
    .B1(addr_i_11_),
    .Y(_07319_)
  );
  sg13g2_a21oi_1 _17114_ (
    .A1(_08310_),
    .A2(_07318_),
    .B1(_07319_),
    .Y(_07320_)
  );
  sg13g2_a21oi_1 _17115_ (
    .A1(_04550_),
    .A2(_01928_),
    .B1(_00064_),
    .Y(_07321_)
  );
  sg13g2_a22oi_1 _17116_ (
    .A1(_03676_),
    .A2(_06331_),
    .B1(_05102_),
    .B2(_07321_),
    .Y(_07322_)
  );
  sg13g2_nand2_1 _17117_ (
    .A(_02141_),
    .B(_06017_),
    .Y(_07323_)
  );
  sg13g2_o21ai_1 _17118_ (
    .A1(addr_i_4_),
    .A2(_07322_),
    .B1(_07323_),
    .Y(_07324_)
  );
  sg13g2_a21oi_1 _17119_ (
    .A1(_00676_),
    .A2(_06331_),
    .B1(_03601_),
    .Y(_07325_)
  );
  sg13g2_a221oi_1 _17120_ (
    .A1(_01537_),
    .A2(_05966_),
    .B1(_06198_),
    .B2(_00664_),
    .C1(addr_i_3_),
    .Y(_07327_)
  );
  sg13g2_a22oi_1 _17121_ (
    .A1(addr_i_3_),
    .A2(_07325_),
    .B1(_07327_),
    .B2(_05302_),
    .Y(_07328_)
  );
  sg13g2_a221oi_1 _17122_ (
    .A1(_05501_),
    .A2(_01923_),
    .B1(_07324_),
    .B2(_02105_),
    .C1(_07328_),
    .Y(_07329_)
  );
  sg13g2_or2_1 _17123_ (
    .A(addr_i_6_),
    .B(_00170_),
    .X(_07330_)
  );
  sg13g2_a221oi_1 _17124_ (
    .A1(_05955_),
    .A2(_07956_),
    .B1(_00768_),
    .B2(_03607_),
    .C1(_00175_),
    .Y(_07331_)
  );
  sg13g2_nor2_1 _17125_ (
    .A(addr_i_6_),
    .B(_07331_),
    .Y(_07332_)
  );
  sg13g2_a221oi_1 _17126_ (
    .A1(_09226_),
    .A2(_06405_),
    .B1(_02514_),
    .B2(_07330_),
    .C1(_07332_),
    .Y(_07333_)
  );
  sg13g2_nand3b_1 _17127_ (
    .A_N(_06441_),
    .B(_01241_),
    .C(addr_i_3_),
    .Y(_07334_)
  );
  sg13g2_o21ai_1 _17128_ (
    .A1(_00873_),
    .A2(_06303_),
    .B1(_07334_),
    .Y(_07335_)
  );
  sg13g2_o21ai_1 _17129_ (
    .A1(addr_i_4_),
    .A2(_02780_),
    .B1(_01911_),
    .Y(_07336_)
  );
  sg13g2_a221oi_1 _17130_ (
    .A1(addr_i_4_),
    .A2(_06021_),
    .B1(_07336_),
    .B2(addr_i_3_),
    .C1(_03270_),
    .Y(_07338_)
  );
  sg13g2_a21o_1 _17131_ (
    .A1(_02343_),
    .A2(_07335_),
    .B1(_07338_),
    .X(_07339_)
  );
  sg13g2_a21oi_1 _17132_ (
    .A1(_07333_),
    .A2(_07339_),
    .B1(_01517_),
    .Y(_07340_)
  );
  sg13g2_a21o_1 _17133_ (
    .A1(_06905_),
    .A2(_07329_),
    .B1(_07340_),
    .X(_07341_)
  );
  sg13g2_o21ai_1 _17134_ (
    .A1(_09348_),
    .A2(_00205_),
    .B1(addr_i_3_),
    .Y(_07342_)
  );
  sg13g2_o21ai_1 _17135_ (
    .A1(_00335_),
    .A2(_02330_),
    .B1(addr_i_4_),
    .Y(_07343_)
  );
  sg13g2_nand3_1 _17136_ (
    .A(_03071_),
    .B(_07342_),
    .C(_07343_),
    .Y(_07344_)
  );
  sg13g2_nor3_1 _17137_ (
    .A(_02304_),
    .B(_03132_),
    .C(_05544_),
    .Y(_07345_)
  );
  sg13g2_nor3_1 _17138_ (
    .A(_04151_),
    .B(_01268_),
    .C(_02179_),
    .Y(_07346_)
  );
  sg13g2_nand2_1 _17139_ (
    .A(_08741_),
    .B(_01539_),
    .Y(_07347_)
  );
  sg13g2_a21oi_1 _17140_ (
    .A1(_04095_),
    .A2(_07347_),
    .B1(_00715_),
    .Y(_07349_)
  );
  sg13g2_or4_1 _17141_ (
    .A(addr_i_9_),
    .B(_07345_),
    .C(_07346_),
    .D(_07349_),
    .X(_07350_)
  );
  sg13g2_nand2_1 _17142_ (
    .A(addr_i_2_),
    .B(_01493_),
    .Y(_07351_)
  );
  sg13g2_nor2_1 _17143_ (
    .A(_00347_),
    .B(_03336_),
    .Y(_07352_)
  );
  sg13g2_o21ai_1 _17144_ (
    .A1(_06501_),
    .A2(_07352_),
    .B1(_00122_),
    .Y(_07353_)
  );
  sg13g2_a21oi_1 _17145_ (
    .A1(_07351_),
    .A2(_07353_),
    .B1(_08674_),
    .Y(_07354_)
  );
  sg13g2_a22oi_1 _17146_ (
    .A1(_01633_),
    .A2(_07344_),
    .B1(_07350_),
    .B2(_07354_),
    .Y(_07355_)
  );
  sg13g2_a22oi_1 _17147_ (
    .A1(addr_i_9_),
    .A2(_07341_),
    .B1(_07355_),
    .B2(addr_i_10_),
    .Y(_07356_)
  );
  sg13g2_nand3_1 _17148_ (
    .A(addr_i_3_),
    .B(addr_i_6_),
    .C(_03424_),
    .Y(_07357_)
  );
  sg13g2_a21oi_1 _17149_ (
    .A1(_02546_),
    .A2(_07357_),
    .B1(addr_i_5_),
    .Y(_07358_)
  );
  sg13g2_o21ai_1 _17150_ (
    .A1(_01962_),
    .A2(_07358_),
    .B1(addr_i_4_),
    .Y(_07360_)
  );
  sg13g2_o21ai_1 _17151_ (
    .A1(_05236_),
    .A2(_03245_),
    .B1(_00400_),
    .Y(_07361_)
  );
  sg13g2_nand3_1 _17152_ (
    .A(_04296_),
    .B(_01343_),
    .C(_07361_),
    .Y(_07362_)
  );
  sg13g2_a22oi_1 _17153_ (
    .A1(_00547_),
    .A2(_00400_),
    .B1(_05021_),
    .B2(addr_i_3_),
    .Y(_07363_)
  );
  sg13g2_a21o_1 _17154_ (
    .A1(_00376_),
    .A2(_01134_),
    .B1(_07363_),
    .X(_07364_)
  );
  sg13g2_nor2_1 _17155_ (
    .A(_00472_),
    .B(_01127_),
    .Y(_07365_)
  );
  sg13g2_o21ai_1 _17156_ (
    .A1(addr_i_4_),
    .A2(_07365_),
    .B1(addr_i_8_),
    .Y(_07366_)
  );
  sg13g2_a221oi_1 _17157_ (
    .A1(addr_i_3_),
    .A2(_07362_),
    .B1(_07364_),
    .B2(addr_i_2_),
    .C1(_07366_),
    .Y(_07367_)
  );
  sg13g2_o21ai_1 _17158_ (
    .A1(_01159_),
    .A2(_01587_),
    .B1(addr_i_3_),
    .Y(_07368_)
  );
  sg13g2_nand3_1 _17159_ (
    .A(_03993_),
    .B(_00007_),
    .C(_02577_),
    .Y(_07369_)
  );
  sg13g2_nand4_1 _17160_ (
    .A(_01520_),
    .B(_00764_),
    .C(_07368_),
    .D(_07369_),
    .Y(_07371_)
  );
  sg13g2_a21oi_1 _17161_ (
    .A1(_01219_),
    .A2(_02553_),
    .B1(addr_i_6_),
    .Y(_07372_)
  );
  sg13g2_a21oi_1 _17162_ (
    .A1(_01368_),
    .A2(_01946_),
    .B1(_03919_),
    .Y(_07373_)
  );
  sg13g2_or4_1 _17163_ (
    .A(_08155_),
    .B(_05590_),
    .C(_07372_),
    .D(_07373_),
    .X(_07374_)
  );
  sg13g2_a22oi_1 _17164_ (
    .A1(_07371_),
    .A2(_07374_),
    .B1(addr_i_8_),
    .B2(_09507_),
    .Y(_07375_)
  );
  sg13g2_a22oi_1 _17165_ (
    .A1(_07360_),
    .A2(_07367_),
    .B1(_00925_),
    .B2(_07375_),
    .Y(_07376_)
  );
  sg13g2_nand3_1 _17166_ (
    .A(addr_i_7_),
    .B(_05648_),
    .C(_04805_),
    .Y(_07377_)
  );
  sg13g2_a21oi_1 _17167_ (
    .A1(_02479_),
    .A2(_02012_),
    .B1(addr_i_3_),
    .Y(_07378_)
  );
  sg13g2_a22oi_1 _17168_ (
    .A1(_01367_),
    .A2(_03853_),
    .B1(_07378_),
    .B2(addr_i_7_),
    .Y(_07379_)
  );
  sg13g2_o21ai_1 _17169_ (
    .A1(_00667_),
    .A2(_04130_),
    .B1(addr_i_6_),
    .Y(_07380_)
  );
  sg13g2_a21oi_1 _17170_ (
    .A1(_07379_),
    .A2(_07380_),
    .B1(addr_i_8_),
    .Y(_07383_)
  );
  sg13g2_o21ai_1 _17171_ (
    .A1(_06715_),
    .A2(_07377_),
    .B1(_07383_),
    .Y(_07384_)
  );
  sg13g2_a21oi_1 _17172_ (
    .A1(_08929_),
    .A2(_06176_),
    .B1(addr_i_5_),
    .Y(_07385_)
  );
  sg13g2_a21oi_1 _17173_ (
    .A1(_00671_),
    .A2(_03915_),
    .B1(_07385_),
    .Y(_07386_)
  );
  sg13g2_o21ai_1 _17174_ (
    .A1(_03139_),
    .A2(_05932_),
    .B1(_00238_),
    .Y(_07387_)
  );
  sg13g2_a21oi_1 _17175_ (
    .A1(_02165_),
    .A2(_07387_),
    .B1(addr_i_7_),
    .Y(_07388_)
  );
  sg13g2_a21oi_1 _17176_ (
    .A1(addr_i_3_),
    .A2(_07386_),
    .B1(_07388_),
    .Y(_07389_)
  );
  sg13g2_a21oi_1 _17177_ (
    .A1(_01672_),
    .A2(_01337_),
    .B1(addr_i_4_),
    .Y(_07390_)
  );
  sg13g2_a21oi_1 _17178_ (
    .A1(_01738_),
    .A2(_04881_),
    .B1(addr_i_5_),
    .Y(_07391_)
  );
  sg13g2_or4_1 _17179_ (
    .A(addr_i_3_),
    .B(_01112_),
    .C(_07390_),
    .D(_07391_),
    .X(_07392_)
  );
  sg13g2_nand4_1 _17180_ (
    .A(addr_i_8_),
    .B(_03340_),
    .C(_07389_),
    .D(_07392_),
    .Y(_07394_)
  );
  sg13g2_a21oi_1 _17181_ (
    .A1(_07384_),
    .A2(_07394_),
    .B1(_01211_),
    .Y(_07395_)
  );
  sg13g2_nor4_1 _17182_ (
    .A(addr_i_11_),
    .B(_07356_),
    .C(_07376_),
    .D(_07395_),
    .Y(_07396_)
  );
  sg13g2_a22oi_1 _17183_ (
    .A1(_07317_),
    .A2(_07320_),
    .B1(_07396_),
    .B2(_00812_),
    .Y(_07397_)
  );
  sg13g2_or2_1 _17184_ (
    .A(_07302_),
    .B(_07397_),
    .X(data_o_30_)
  );
  sg13g2_a21oi_1 _17185_ (
    .A1(_08431_),
    .A2(_01290_),
    .B1(_02136_),
    .Y(_07398_)
  );
  sg13g2_a22oi_1 _17186_ (
    .A1(addr_i_4_),
    .A2(_07480_),
    .B1(_03980_),
    .B2(addr_i_7_),
    .Y(_07399_)
  );
  sg13g2_o21ai_1 _17187_ (
    .A1(_00302_),
    .A2(_01049_),
    .B1(addr_i_3_),
    .Y(_07400_)
  );
  sg13g2_nor4_1 _17188_ (
    .A(_04483_),
    .B(_02265_),
    .C(_01402_),
    .D(_02069_),
    .Y(_07401_)
  );
  sg13g2_nor2_1 _17189_ (
    .A(_04815_),
    .B(_05883_),
    .Y(_07402_)
  );
  sg13g2_nand4_1 _17190_ (
    .A(_02530_),
    .B(_08232_),
    .C(_07401_),
    .D(_07402_),
    .Y(_07404_)
  );
  sg13g2_o21ai_1 _17191_ (
    .A1(_07399_),
    .A2(_07400_),
    .B1(_07404_),
    .Y(_07405_)
  );
  sg13g2_o21ai_1 _17192_ (
    .A1(_07398_),
    .A2(_07405_),
    .B1(addr_i_8_),
    .Y(_07406_)
  );
  sg13g2_o21ai_1 _17193_ (
    .A1(_06795_),
    .A2(_06806_),
    .B1(addr_i_3_),
    .Y(_07407_)
  );
  sg13g2_o21ai_1 _17194_ (
    .A1(_05501_),
    .A2(_07647_),
    .B1(_01653_),
    .Y(_07408_)
  );
  sg13g2_nand3_1 _17195_ (
    .A(_02467_),
    .B(_07407_),
    .C(_07408_),
    .Y(_07409_)
  );
  sg13g2_o21ai_1 _17196_ (
    .A1(_05258_),
    .A2(_00333_),
    .B1(_00749_),
    .Y(_07410_)
  );
  sg13g2_a21oi_1 _17197_ (
    .A1(_00731_),
    .A2(_00547_),
    .B1(_00445_),
    .Y(_07411_)
  );
  sg13g2_a22oi_1 _17198_ (
    .A1(_00778_),
    .A2(_07410_),
    .B1(_07411_),
    .B2(_04915_),
    .Y(_07412_)
  );
  sg13g2_nand2_1 _17199_ (
    .A(_00145_),
    .B(_02569_),
    .Y(_07413_)
  );
  sg13g2_a22oi_1 _17200_ (
    .A1(_03348_),
    .A2(_07413_),
    .B1(addr_i_4_),
    .B2(_02772_),
    .Y(_07415_)
  );
  sg13g2_a21oi_1 _17201_ (
    .A1(addr_i_4_),
    .A2(_07412_),
    .B1(_07415_),
    .Y(_07416_)
  );
  sg13g2_a22oi_1 _17202_ (
    .A1(addr_i_7_),
    .A2(_07409_),
    .B1(_07416_),
    .B2(addr_i_8_),
    .Y(_07417_)
  );
  sg13g2_nor2_1 _17203_ (
    .A(_01452_),
    .B(_07417_),
    .Y(_07418_)
  );
  sg13g2_nand3_1 _17204_ (
    .A(_00339_),
    .B(_02656_),
    .C(_03871_),
    .Y(_07419_)
  );
  sg13g2_o21ai_1 _17205_ (
    .A1(_08885_),
    .A2(_03194_),
    .B1(addr_i_3_),
    .Y(_07420_)
  );
  sg13g2_a21oi_1 _17206_ (
    .A1(_00849_),
    .A2(_07420_),
    .B1(_00230_),
    .Y(_07421_)
  );
  sg13g2_a221oi_1 _17207_ (
    .A1(_05081_),
    .A2(_00783_),
    .B1(_04754_),
    .B2(_09497_),
    .C1(_00746_),
    .Y(_07422_)
  );
  sg13g2_o21ai_1 _17208_ (
    .A1(_02203_),
    .A2(_02161_),
    .B1(addr_i_2_),
    .Y(_07423_)
  );
  sg13g2_a21oi_1 _17209_ (
    .A1(_07422_),
    .A2(_07423_),
    .B1(_06905_),
    .Y(_07424_)
  );
  sg13g2_a22oi_1 _17210_ (
    .A1(_09487_),
    .A2(_07419_),
    .B1(_07421_),
    .B2(_07424_),
    .Y(_07426_)
  );
  sg13g2_nor2_1 _17211_ (
    .A(_00492_),
    .B(_01480_),
    .Y(_07427_)
  );
  sg13g2_nor3_1 _17212_ (
    .A(addr_i_2_),
    .B(_00372_),
    .C(_02389_),
    .Y(_07428_)
  );
  sg13g2_o21ai_1 _17213_ (
    .A1(addr_i_3_),
    .A2(_05651_),
    .B1(_02708_),
    .Y(_07429_)
  );
  sg13g2_o21ai_1 _17214_ (
    .A1(_02287_),
    .A2(_07429_),
    .B1(addr_i_7_),
    .Y(_07430_)
  );
  sg13g2_a22oi_1 _17215_ (
    .A1(addr_i_4_),
    .A2(_02755_),
    .B1(_01107_),
    .B2(addr_i_3_),
    .Y(_07431_)
  );
  sg13g2_o21ai_1 _17216_ (
    .A1(_02922_),
    .A2(_07431_),
    .B1(_01878_),
    .Y(_07432_)
  );
  sg13g2_o21ai_1 _17217_ (
    .A1(_07428_),
    .A2(_07430_),
    .B1(_07432_),
    .Y(_07433_)
  );
  sg13g2_a22oi_1 _17218_ (
    .A1(_02948_),
    .A2(_07427_),
    .B1(_07433_),
    .B2(addr_i_8_),
    .Y(_07434_)
  );
  sg13g2_a22oi_1 _17219_ (
    .A1(addr_i_8_),
    .A2(_07426_),
    .B1(_07434_),
    .B2(_02221_),
    .Y(_07435_)
  );
  sg13g2_a21oi_1 _17220_ (
    .A1(addr_i_6_),
    .A2(_00090_),
    .B1(_06541_),
    .Y(_07437_)
  );
  sg13g2_a21oi_1 _17221_ (
    .A1(_02623_),
    .A2(_00583_),
    .B1(_01424_),
    .Y(_07438_)
  );
  sg13g2_o21ai_1 _17222_ (
    .A1(addr_i_3_),
    .A2(_07437_),
    .B1(_07438_),
    .Y(_07439_)
  );
  sg13g2_o21ai_1 _17223_ (
    .A1(_02639_),
    .A2(_02641_),
    .B1(addr_i_5_),
    .Y(_07440_)
  );
  sg13g2_o21ai_1 _17224_ (
    .A1(_00716_),
    .A2(_02437_),
    .B1(_07440_),
    .Y(_07441_)
  );
  sg13g2_o21ai_1 _17225_ (
    .A1(_02437_),
    .A2(_04095_),
    .B1(addr_i_8_),
    .Y(_07442_)
  );
  sg13g2_a221oi_1 _17226_ (
    .A1(addr_i_4_),
    .A2(_07439_),
    .B1(_07441_),
    .B2(addr_i_2_),
    .C1(_07442_),
    .Y(_07443_)
  );
  sg13g2_nand2b_1 _17227_ (
    .A_N(_07443_),
    .B(_00773_),
    .Y(_07444_)
  );
  sg13g2_o21ai_1 _17228_ (
    .A1(_02215_),
    .A2(_03812_),
    .B1(addr_i_2_),
    .Y(_07445_)
  );
  sg13g2_o21ai_1 _17229_ (
    .A1(_00961_),
    .A2(_06473_),
    .B1(_07445_),
    .Y(_07446_)
  );
  sg13g2_a21oi_1 _17230_ (
    .A1(_02815_),
    .A2(_02529_),
    .B1(addr_i_3_),
    .Y(_07448_)
  );
  sg13g2_o21ai_1 _17231_ (
    .A1(_00597_),
    .A2(_07448_),
    .B1(_01517_),
    .Y(_07449_)
  );
  sg13g2_a21oi_1 _17232_ (
    .A1(_00021_),
    .A2(_00434_),
    .B1(_00522_),
    .Y(_07450_)
  );
  sg13g2_o21ai_1 _17233_ (
    .A1(_04400_),
    .A2(_07450_),
    .B1(addr_i_5_),
    .Y(_07451_)
  );
  sg13g2_nand2_1 _17234_ (
    .A(_07449_),
    .B(_07451_),
    .Y(_07452_)
  );
  sg13g2_a22oi_1 _17235_ (
    .A1(addr_i_4_),
    .A2(_07446_),
    .B1(_07452_),
    .B2(addr_i_8_),
    .Y(_07453_)
  );
  sg13g2_a21oi_1 _17236_ (
    .A1(_05036_),
    .A2(_02020_),
    .B1(addr_i_4_),
    .Y(_07454_)
  );
  sg13g2_a21oi_1 _17237_ (
    .A1(addr_i_4_),
    .A2(_06473_),
    .B1(_07454_),
    .Y(_07455_)
  );
  sg13g2_o21ai_1 _17238_ (
    .A1(_01674_),
    .A2(_07455_),
    .B1(_00831_),
    .Y(_07456_)
  );
  sg13g2_nand3_1 _17239_ (
    .A(_01834_),
    .B(_03324_),
    .C(_07420_),
    .Y(_07457_)
  );
  sg13g2_o21ai_1 _17240_ (
    .A1(_01155_),
    .A2(_07457_),
    .B1(addr_i_8_),
    .Y(_07459_)
  );
  sg13g2_a221oi_1 _17241_ (
    .A1(_01662_),
    .A2(_02839_),
    .B1(_07456_),
    .B2(addr_i_7_),
    .C1(_07459_),
    .Y(_07460_)
  );
  sg13g2_nand2_1 _17242_ (
    .A(_07779_),
    .B(_04769_),
    .Y(_07461_)
  );
  sg13g2_o21ai_1 _17243_ (
    .A1(addr_i_4_),
    .A2(_03288_),
    .B1(_07713_),
    .Y(_07462_)
  );
  sg13g2_a22oi_1 _17244_ (
    .A1(_00145_),
    .A2(_07461_),
    .B1(_07462_),
    .B2(_03820_),
    .Y(_07463_)
  );
  sg13g2_a21oi_1 _17245_ (
    .A1(_02602_),
    .A2(_00333_),
    .B1(_02343_),
    .Y(_07464_)
  );
  sg13g2_nand3_1 _17246_ (
    .A(_05281_),
    .B(_01373_),
    .C(_01976_),
    .Y(_07465_)
  );
  sg13g2_a21oi_1 _17247_ (
    .A1(_06552_),
    .A2(_07465_),
    .B1(_04108_),
    .Y(_07466_)
  );
  sg13g2_nor4_1 _17248_ (
    .A(addr_i_7_),
    .B(_00472_),
    .C(_07464_),
    .D(_07466_),
    .Y(_07467_)
  );
  sg13g2_or3_1 _17249_ (
    .A(addr_i_8_),
    .B(_07463_),
    .C(_07467_),
    .X(_07468_)
  );
  sg13g2_nand3b_1 _17250_ (
    .A_N(_07460_),
    .B(_07468_),
    .C(_01174_),
    .Y(_07470_)
  );
  sg13g2_o21ai_1 _17251_ (
    .A1(_07444_),
    .A2(_07453_),
    .B1(_07470_),
    .Y(_07471_)
  );
  sg13g2_a22oi_1 _17252_ (
    .A1(_07406_),
    .A2(_07418_),
    .B1(_07435_),
    .B2(_07471_),
    .Y(_07472_)
  );
  sg13g2_o21ai_1 _17253_ (
    .A1(_05524_),
    .A2(_01014_),
    .B1(_08696_),
    .Y(_07473_)
  );
  sg13g2_a21oi_1 _17254_ (
    .A1(_01588_),
    .A2(_07473_),
    .B1(addr_i_7_),
    .Y(_07474_)
  );
  sg13g2_nor3_1 _17255_ (
    .A(_08696_),
    .B(_08144_),
    .C(_00247_),
    .Y(_07475_)
  );
  sg13g2_a22oi_1 _17256_ (
    .A1(_00445_),
    .A2(_09509_),
    .B1(_07475_),
    .B2(_06375_),
    .Y(_07476_)
  );
  sg13g2_o21ai_1 _17257_ (
    .A1(_07474_),
    .A2(_07476_),
    .B1(addr_i_3_),
    .Y(_07477_)
  );
  sg13g2_o21ai_1 _17258_ (
    .A1(_02213_),
    .A2(_07248_),
    .B1(_03226_),
    .Y(_07478_)
  );
  sg13g2_a21oi_1 _17259_ (
    .A1(_01354_),
    .A2(_00131_),
    .B1(_00778_),
    .Y(_07479_)
  );
  sg13g2_a22oi_1 _17260_ (
    .A1(_07824_),
    .A2(_07478_),
    .B1(_07479_),
    .B2(addr_i_8_),
    .Y(_07481_)
  );
  sg13g2_nand2_1 _17261_ (
    .A(_04068_),
    .B(_00801_),
    .Y(_07482_)
  );
  sg13g2_o21ai_1 _17262_ (
    .A1(_06398_),
    .A2(_00334_),
    .B1(_01215_),
    .Y(_07483_)
  );
  sg13g2_a21oi_1 _17263_ (
    .A1(_04671_),
    .A2(_07483_),
    .B1(addr_i_7_),
    .Y(_07484_)
  );
  sg13g2_a22oi_1 _17264_ (
    .A1(addr_i_4_),
    .A2(_07482_),
    .B1(_07484_),
    .B2(_06695_),
    .Y(_07485_)
  );
  sg13g2_a22oi_1 _17265_ (
    .A1(_07477_),
    .A2(_07481_),
    .B1(addr_i_9_),
    .B2(_07485_),
    .Y(_07486_)
  );
  sg13g2_o21ai_1 _17266_ (
    .A1(_03886_),
    .A2(_03494_),
    .B1(addr_i_10_),
    .Y(_07487_)
  );
  sg13g2_o21ai_1 _17267_ (
    .A1(_02399_),
    .A2(_07486_),
    .B1(_07487_),
    .Y(_07488_)
  );
  sg13g2_and2_1 _17268_ (
    .A(addr_i_11_),
    .B(_07488_),
    .X(_07489_)
  );
  sg13g2_a21oi_1 _17269_ (
    .A1(_03051_),
    .A2(_07472_),
    .B1(_07489_),
    .Y(_07490_)
  );
  sg13g2_a22oi_1 _17270_ (
    .A1(_03288_),
    .A2(_01830_),
    .B1(_00205_),
    .B2(_01011_),
    .Y(_07493_)
  );
  sg13g2_xnor2_1 _17271_ (
    .A(_03709_),
    .B(_00583_),
    .Y(_07494_)
  );
  sg13g2_a21oi_1 _17272_ (
    .A1(_06386_),
    .A2(_06851_),
    .B1(_00718_),
    .Y(_07495_)
  );
  sg13g2_a221oi_1 _17273_ (
    .A1(_00586_),
    .A2(_01033_),
    .B1(_07494_),
    .B2(_00199_),
    .C1(_07495_),
    .Y(_07496_)
  );
  sg13g2_nor2_1 _17274_ (
    .A(_01274_),
    .B(_07496_),
    .Y(_07497_)
  );
  sg13g2_a22oi_1 _17275_ (
    .A1(_03582_),
    .A2(_07493_),
    .B1(_07497_),
    .B2(_00374_),
    .Y(_07498_)
  );
  sg13g2_nand2_1 _17276_ (
    .A(_05236_),
    .B(_00319_),
    .Y(_07499_)
  );
  sg13g2_nand3_1 _17277_ (
    .A(addr_i_3_),
    .B(_04429_),
    .C(_05910_),
    .Y(_07500_)
  );
  sg13g2_a21oi_1 _17278_ (
    .A1(_07499_),
    .A2(_07500_),
    .B1(_00145_),
    .Y(_07501_)
  );
  sg13g2_o21ai_1 _17279_ (
    .A1(addr_i_7_),
    .A2(_01472_),
    .B1(_02462_),
    .Y(_07502_)
  );
  sg13g2_nand2_1 _17280_ (
    .A(_01544_),
    .B(_07502_),
    .Y(_07504_)
  );
  sg13g2_o21ai_1 _17281_ (
    .A1(_07501_),
    .A2(_07504_),
    .B1(addr_i_5_),
    .Y(_07505_)
  );
  sg13g2_a21oi_1 _17282_ (
    .A1(_08929_),
    .A2(_00210_),
    .B1(_01567_),
    .Y(_07506_)
  );
  sg13g2_o21ai_1 _17283_ (
    .A1(_09513_),
    .A2(_04399_),
    .B1(_07506_),
    .Y(_07507_)
  );
  sg13g2_nor2_1 _17284_ (
    .A(_01948_),
    .B(_00522_),
    .Y(_07508_)
  );
  sg13g2_a21oi_1 _17285_ (
    .A1(_00949_),
    .A2(_07507_),
    .B1(_07508_),
    .Y(_07509_)
  );
  sg13g2_nand3_1 _17286_ (
    .A(_07498_),
    .B(_07505_),
    .C(_07509_),
    .Y(_07510_)
  );
  sg13g2_a21oi_1 _17287_ (
    .A1(addr_i_4_),
    .A2(_00702_),
    .B1(_02108_),
    .Y(_07511_)
  );
  sg13g2_o21ai_1 _17288_ (
    .A1(_05346_),
    .A2(_00308_),
    .B1(addr_i_6_),
    .Y(_07512_)
  );
  sg13g2_o21ai_1 _17289_ (
    .A1(_00463_),
    .A2(_07511_),
    .B1(_07512_),
    .Y(_07513_)
  );
  sg13g2_a21oi_1 _17290_ (
    .A1(_01976_),
    .A2(_02207_),
    .B1(_00342_),
    .Y(_07515_)
  );
  sg13g2_nor4_1 _17291_ (
    .A(_00934_),
    .B(_01274_),
    .C(_01869_),
    .D(_07515_),
    .Y(_07516_)
  );
  sg13g2_o21ai_1 _17292_ (
    .A1(_01659_),
    .A2(_02441_),
    .B1(_00479_),
    .Y(_07517_)
  );
  sg13g2_a221oi_1 _17293_ (
    .A1(_01310_),
    .A2(_07513_),
    .B1(_07516_),
    .B2(_07517_),
    .C1(addr_i_9_),
    .Y(_07518_)
  );
  sg13g2_o21ai_1 _17294_ (
    .A1(_05590_),
    .A2(_04316_),
    .B1(addr_i_2_),
    .Y(_07519_)
  );
  sg13g2_a21oi_1 _17295_ (
    .A1(_04119_),
    .A2(_02405_),
    .B1(_01229_),
    .Y(_07520_)
  );
  sg13g2_a21oi_1 _17296_ (
    .A1(_07519_),
    .A2(_07520_),
    .B1(addr_i_4_),
    .Y(_07521_)
  );
  sg13g2_a22oi_1 _17297_ (
    .A1(_01580_),
    .A2(_03112_),
    .B1(_05588_),
    .B2(_07521_),
    .Y(_07522_)
  );
  sg13g2_a21oi_1 _17298_ (
    .A1(_00299_),
    .A2(_04330_),
    .B1(_08000_),
    .Y(_07523_)
  );
  sg13g2_o21ai_1 _17299_ (
    .A1(addr_i_2_),
    .A2(_06693_),
    .B1(_05599_),
    .Y(_07524_)
  );
  sg13g2_o21ai_1 _17300_ (
    .A1(_07523_),
    .A2(_07524_),
    .B1(addr_i_4_),
    .Y(_07526_)
  );
  sg13g2_nand3_1 _17301_ (
    .A(_07518_),
    .B(_07522_),
    .C(_07526_),
    .Y(_07527_)
  );
  sg13g2_o21ai_1 _17302_ (
    .A1(_07498_),
    .A2(_07518_),
    .B1(addr_i_8_),
    .Y(_07528_)
  );
  sg13g2_nand3_1 _17303_ (
    .A(_07510_),
    .B(_07527_),
    .C(_07528_),
    .Y(_07529_)
  );
  sg13g2_nand3_1 _17304_ (
    .A(addr_i_6_),
    .B(_00994_),
    .C(_01087_),
    .Y(_07530_)
  );
  sg13g2_o21ai_1 _17305_ (
    .A1(addr_i_5_),
    .A2(_07061_),
    .B1(addr_i_4_),
    .Y(_07531_)
  );
  sg13g2_nand4_1 _17306_ (
    .A(_00484_),
    .B(_03413_),
    .C(_05689_),
    .D(_07531_),
    .Y(_07532_)
  );
  sg13g2_nand3_1 _17307_ (
    .A(addr_i_3_),
    .B(_07530_),
    .C(_07532_),
    .Y(_07533_)
  );
  sg13g2_nor2_1 _17308_ (
    .A(addr_i_7_),
    .B(_05379_),
    .Y(_07534_)
  );
  sg13g2_a21o_1 _17309_ (
    .A1(_05324_),
    .A2(_02166_),
    .B1(_07534_),
    .X(_07535_)
  );
  sg13g2_a21oi_1 _17310_ (
    .A1(_00050_),
    .A2(_02440_),
    .B1(addr_i_3_),
    .Y(_07537_)
  );
  sg13g2_a22oi_1 _17311_ (
    .A1(_00648_),
    .A2(_07535_),
    .B1(_07537_),
    .B2(_02420_),
    .Y(_07538_)
  );
  sg13g2_nand2_1 _17312_ (
    .A(_07533_),
    .B(_07538_),
    .Y(_07539_)
  );
  sg13g2_o21ai_1 _17313_ (
    .A1(_07636_),
    .A2(_03012_),
    .B1(addr_i_4_),
    .Y(_07540_)
  );
  sg13g2_o21ai_1 _17314_ (
    .A1(_04086_),
    .A2(_09083_),
    .B1(_05379_),
    .Y(_07541_)
  );
  sg13g2_o21ai_1 _17315_ (
    .A1(_06530_),
    .A2(_06541_),
    .B1(_00535_),
    .Y(_07542_)
  );
  sg13g2_nand3_1 _17316_ (
    .A(_07540_),
    .B(_07541_),
    .C(_07542_),
    .Y(_07543_)
  );
  sg13g2_nor2_1 _17317_ (
    .A(_04804_),
    .B(_02722_),
    .Y(_07544_)
  );
  sg13g2_a21oi_1 _17318_ (
    .A1(_02086_),
    .A2(_03289_),
    .B1(_07544_),
    .Y(_07545_)
  );
  sg13g2_o21ai_1 _17319_ (
    .A1(_00260_),
    .A2(_02369_),
    .B1(_03523_),
    .Y(_07546_)
  );
  sg13g2_o21ai_1 _17320_ (
    .A1(_00665_),
    .A2(_07545_),
    .B1(_07546_),
    .Y(_07548_)
  );
  sg13g2_a22oi_1 _17321_ (
    .A1(addr_i_7_),
    .A2(_07543_),
    .B1(_07548_),
    .B2(addr_i_8_),
    .Y(_07549_)
  );
  sg13g2_a22oi_1 _17322_ (
    .A1(addr_i_8_),
    .A2(_07539_),
    .B1(_07549_),
    .B2(_00385_),
    .Y(_07550_)
  );
  sg13g2_a21o_1 _17323_ (
    .A1(addr_i_4_),
    .A2(_06790_),
    .B1(_00119_),
    .X(_07551_)
  );
  sg13g2_a21oi_1 _17324_ (
    .A1(_00739_),
    .A2(_02032_),
    .B1(addr_i_4_),
    .Y(_07552_)
  );
  sg13g2_a21oi_1 _17325_ (
    .A1(addr_i_3_),
    .A2(_07551_),
    .B1(_07552_),
    .Y(_07553_)
  );
  sg13g2_nor2_1 _17326_ (
    .A(_02733_),
    .B(_08796_),
    .Y(_07554_)
  );
  sg13g2_nor2_1 _17327_ (
    .A(_07554_),
    .B(_02330_),
    .Y(_07555_)
  );
  sg13g2_o21ai_1 _17328_ (
    .A1(_01086_),
    .A2(_01910_),
    .B1(_01970_),
    .Y(_07556_)
  );
  sg13g2_nand2_1 _17329_ (
    .A(_00484_),
    .B(_02218_),
    .Y(_07557_)
  );
  sg13g2_a21oi_1 _17330_ (
    .A1(_04539_),
    .A2(_07557_),
    .B1(_02535_),
    .Y(_07559_)
  );
  sg13g2_nand4_1 _17331_ (
    .A(_07555_),
    .B(_05864_),
    .C(_07556_),
    .D(_07559_),
    .Y(_07560_)
  );
  sg13g2_o21ai_1 _17332_ (
    .A1(_03494_),
    .A2(_07553_),
    .B1(_07560_),
    .Y(_07561_)
  );
  sg13g2_o21ai_1 _17333_ (
    .A1(_00637_),
    .A2(_04937_),
    .B1(_00199_),
    .Y(_07562_)
  );
  sg13g2_a21oi_1 _17334_ (
    .A1(_00878_),
    .A2(_07562_),
    .B1(addr_i_7_),
    .Y(_07563_)
  );
  sg13g2_a21oi_1 _17335_ (
    .A1(_00566_),
    .A2(_03405_),
    .B1(_00744_),
    .Y(_07564_)
  );
  sg13g2_or2_1 _17336_ (
    .A(_07563_),
    .B(_07564_),
    .X(_07565_)
  );
  sg13g2_a21oi_1 _17337_ (
    .A1(_03540_),
    .A2(_01077_),
    .B1(_00381_),
    .Y(_07566_)
  );
  sg13g2_a21oi_1 _17338_ (
    .A1(addr_i_7_),
    .A2(_01160_),
    .B1(addr_i_5_),
    .Y(_07567_)
  );
  sg13g2_nor4_1 _17339_ (
    .A(addr_i_3_),
    .B(_00257_),
    .C(_07566_),
    .D(_07567_),
    .Y(_07568_)
  );
  sg13g2_nor2_1 _17340_ (
    .A(addr_i_7_),
    .B(_01459_),
    .Y(_07570_)
  );
  sg13g2_o21ai_1 _17341_ (
    .A1(_00695_),
    .A2(_07570_),
    .B1(_02604_),
    .Y(_07571_)
  );
  sg13g2_a22oi_1 _17342_ (
    .A1(addr_i_3_),
    .A2(_07565_),
    .B1(_07568_),
    .B2(_07571_),
    .Y(_07572_)
  );
  sg13g2_nor4_1 _17343_ (
    .A(addr_i_10_),
    .B(_07550_),
    .C(_07561_),
    .D(_07572_),
    .Y(_07573_)
  );
  sg13g2_a21o_1 _17344_ (
    .A1(addr_i_10_),
    .A2(_07529_),
    .B1(_07573_),
    .X(_07574_)
  );
  sg13g2_nand3b_1 _17345_ (
    .A_N(_02198_),
    .B(addr_i_4_),
    .C(_01791_),
    .Y(_07575_)
  );
  sg13g2_nand3_1 _17346_ (
    .A(_00554_),
    .B(_02471_),
    .C(_00404_),
    .Y(_07576_)
  );
  sg13g2_a21oi_1 _17347_ (
    .A1(addr_i_4_),
    .A2(_02471_),
    .B1(_00155_),
    .Y(_07577_)
  );
  sg13g2_a21oi_1 _17348_ (
    .A1(_07575_),
    .A2(_07576_),
    .B1(_07577_),
    .Y(_07578_)
  );
  sg13g2_nor2_1 _17349_ (
    .A(_04782_),
    .B(_00946_),
    .Y(_07579_)
  );
  sg13g2_a22oi_1 _17350_ (
    .A1(addr_i_2_),
    .A2(_05231_),
    .B1(_00096_),
    .B2(_00354_),
    .Y(_07581_)
  );
  sg13g2_a22oi_1 _17351_ (
    .A1(_00554_),
    .A2(_07579_),
    .B1(_07581_),
    .B2(_02105_),
    .Y(_07582_)
  );
  sg13g2_nor2_1 _17352_ (
    .A(_05546_),
    .B(_00679_),
    .Y(_07583_)
  );
  sg13g2_nor3_1 _17353_ (
    .A(_02542_),
    .B(_07582_),
    .C(_07583_),
    .Y(_07584_)
  );
  sg13g2_o21ai_1 _17354_ (
    .A1(addr_i_3_),
    .A2(_07578_),
    .B1(_07584_),
    .Y(_07585_)
  );
  sg13g2_nor3_1 _17355_ (
    .A(addr_i_3_),
    .B(_00014_),
    .C(_06264_),
    .Y(_07586_)
  );
  sg13g2_or2_1 _17356_ (
    .A(_01275_),
    .B(_07586_),
    .X(_07587_)
  );
  sg13g2_nand2_1 _17357_ (
    .A(_05357_),
    .B(_05021_),
    .Y(_07588_)
  );
  sg13g2_a221oi_1 _17358_ (
    .A1(addr_i_3_),
    .A2(_06663_),
    .B1(_07587_),
    .B2(_07588_),
    .C1(_02535_),
    .Y(_07589_)
  );
  sg13g2_nand2_1 _17359_ (
    .A(_03431_),
    .B(_00422_),
    .Y(_07590_)
  );
  sg13g2_a22oi_1 _17360_ (
    .A1(addr_i_3_),
    .A2(_03323_),
    .B1(_07590_),
    .B2(_01481_),
    .Y(_07592_)
  );
  sg13g2_a22oi_1 _17361_ (
    .A1(_02604_),
    .A2(_07585_),
    .B1(_07589_),
    .B2(_07592_),
    .Y(_07593_)
  );
  sg13g2_a21oi_1 _17362_ (
    .A1(_00381_),
    .A2(_04095_),
    .B1(addr_i_2_),
    .Y(_07594_)
  );
  sg13g2_inv_1 _17363_ (
    .A(_02179_),
    .Y(_07595_)
  );
  sg13g2_o21ai_1 _17364_ (
    .A1(_02792_),
    .A2(_07594_),
    .B1(_07595_),
    .Y(_07596_)
  );
  sg13g2_nand3_1 _17365_ (
    .A(addr_i_4_),
    .B(_07326_),
    .C(_09393_),
    .Y(_07597_)
  );
  sg13g2_nand3_1 _17366_ (
    .A(_05125_),
    .B(_01168_),
    .C(_07597_),
    .Y(_07598_)
  );
  sg13g2_a21oi_1 _17367_ (
    .A1(_04618_),
    .A2(_04371_),
    .B1(_01494_),
    .Y(_07599_)
  );
  sg13g2_nand2_1 _17368_ (
    .A(_07598_),
    .B(_07599_),
    .Y(_07600_)
  );
  sg13g2_a21oi_1 _17369_ (
    .A1(_01757_),
    .A2(_01768_),
    .B1(addr_i_3_),
    .Y(_07601_)
  );
  sg13g2_a21oi_1 _17370_ (
    .A1(addr_i_3_),
    .A2(_07480_),
    .B1(_07601_),
    .Y(_07604_)
  );
  sg13g2_nor2_1 _17371_ (
    .A(_04373_),
    .B(_07604_),
    .Y(_07605_)
  );
  sg13g2_a21oi_1 _17372_ (
    .A1(_07569_),
    .A2(_01182_),
    .B1(addr_i_6_),
    .Y(_07606_)
  );
  sg13g2_o21ai_1 _17373_ (
    .A1(_07605_),
    .A2(_07606_),
    .B1(_01666_),
    .Y(_07607_)
  );
  sg13g2_nand3_1 _17374_ (
    .A(_07596_),
    .B(_07600_),
    .C(_07607_),
    .Y(_07608_)
  );
  sg13g2_nand2_1 _17375_ (
    .A(_00320_),
    .B(_06052_),
    .Y(_07609_)
  );
  sg13g2_a21o_1 _17376_ (
    .A1(_02799_),
    .A2(_04114_),
    .B1(_02086_),
    .X(_07610_)
  );
  sg13g2_a21oi_1 _17377_ (
    .A1(_03478_),
    .A2(_07610_),
    .B1(addr_i_7_),
    .Y(_07611_)
  );
  sg13g2_a22oi_1 _17378_ (
    .A1(_00262_),
    .A2(_07609_),
    .B1(_07611_),
    .B2(_01286_),
    .Y(_07612_)
  );
  sg13g2_nor2_1 _17379_ (
    .A(addr_i_8_),
    .B(_07612_),
    .Y(_07613_)
  );
  sg13g2_o21ai_1 _17380_ (
    .A1(_07608_),
    .A2(_07613_),
    .B1(addr_i_9_),
    .Y(_07615_)
  );
  sg13g2_a21o_1 _17381_ (
    .A1(_07593_),
    .A2(_07615_),
    .B1(addr_i_10_),
    .X(_07616_)
  );
  sg13g2_a21oi_1 _17382_ (
    .A1(addr_i_3_),
    .A2(_02437_),
    .B1(_05025_),
    .Y(_07617_)
  );
  sg13g2_o21ai_1 _17383_ (
    .A1(_00838_),
    .A2(_00338_),
    .B1(_00645_),
    .Y(_07618_)
  );
  sg13g2_o21ai_1 _17384_ (
    .A1(_02755_),
    .A2(_07617_),
    .B1(_07618_),
    .Y(_07619_)
  );
  sg13g2_o21ai_1 _17385_ (
    .A1(_01194_),
    .A2(_00017_),
    .B1(addr_i_3_),
    .Y(_07620_)
  );
  sg13g2_a22oi_1 _17386_ (
    .A1(_06054_),
    .A2(_04483_),
    .B1(_01977_),
    .B2(_01577_),
    .Y(_07621_)
  );
  sg13g2_a21oi_1 _17387_ (
    .A1(_07620_),
    .A2(_07621_),
    .B1(addr_i_6_),
    .Y(_07622_)
  );
  sg13g2_nor3_1 _17388_ (
    .A(_00113_),
    .B(_07619_),
    .C(_07622_),
    .Y(_07623_)
  );
  sg13g2_nand2_1 _17389_ (
    .A(_04218_),
    .B(_01680_),
    .Y(_07624_)
  );
  sg13g2_nand3_1 _17390_ (
    .A(_04396_),
    .B(_00427_),
    .C(_07624_),
    .Y(_07626_)
  );
  sg13g2_nand2_1 _17391_ (
    .A(_08155_),
    .B(_03721_),
    .Y(_07627_)
  );
  sg13g2_o21ai_1 _17392_ (
    .A1(_08299_),
    .A2(_02626_),
    .B1(_05025_),
    .Y(_07628_)
  );
  sg13g2_nand3_1 _17393_ (
    .A(_00618_),
    .B(_07627_),
    .C(_07628_),
    .Y(_07629_)
  );
  sg13g2_o21ai_1 _17394_ (
    .A1(_03914_),
    .A2(_07001_),
    .B1(_00666_),
    .Y(_07630_)
  );
  sg13g2_nand2_1 _17395_ (
    .A(_03617_),
    .B(_07630_),
    .Y(_07631_)
  );
  sg13g2_a221oi_1 _17396_ (
    .A1(addr_i_5_),
    .A2(_07626_),
    .B1(_07629_),
    .B2(addr_i_3_),
    .C1(_07631_),
    .Y(_07632_)
  );
  sg13g2_o21ai_1 _17397_ (
    .A1(_00569_),
    .A2(_02792_),
    .B1(_03292_),
    .Y(_07633_)
  );
  sg13g2_a21oi_1 _17398_ (
    .A1(addr_i_3_),
    .A2(_01483_),
    .B1(_08045_),
    .Y(_07634_)
  );
  sg13g2_nand2_1 _17399_ (
    .A(_07633_),
    .B(_07634_),
    .Y(_07635_)
  );
  sg13g2_o21ai_1 _17400_ (
    .A1(_07623_),
    .A2(_07632_),
    .B1(_07635_),
    .Y(_07637_)
  );
  sg13g2_a21oi_1 _17401_ (
    .A1(_01004_),
    .A2(_02254_),
    .B1(addr_i_3_),
    .Y(_07638_)
  );
  sg13g2_a21oi_1 _17402_ (
    .A1(_01508_),
    .A2(_00268_),
    .B1(_07638_),
    .Y(_07639_)
  );
  sg13g2_nor2_1 _17403_ (
    .A(addr_i_6_),
    .B(_07639_),
    .Y(_07640_)
  );
  sg13g2_nand2_1 _17404_ (
    .A(_04384_),
    .B(_08221_),
    .Y(_07641_)
  );
  sg13g2_a221oi_1 _17405_ (
    .A1(_05833_),
    .A2(_00448_),
    .B1(_07641_),
    .B2(addr_i_4_),
    .C1(_05883_),
    .Y(_07642_)
  );
  sg13g2_a21oi_1 _17406_ (
    .A1(addr_i_3_),
    .A2(_05457_),
    .B1(_08144_),
    .Y(_07643_)
  );
  sg13g2_o21ai_1 _17407_ (
    .A1(addr_i_4_),
    .A2(_01437_),
    .B1(_00052_),
    .Y(_07644_)
  );
  sg13g2_a221oi_1 _17408_ (
    .A1(_00029_),
    .A2(_07643_),
    .B1(_07644_),
    .B2(_03993_),
    .C1(_03849_),
    .Y(_07645_)
  );
  sg13g2_o21ai_1 _17409_ (
    .A1(_02530_),
    .A2(_07642_),
    .B1(_07645_),
    .Y(_07646_)
  );
  sg13g2_o21ai_1 _17410_ (
    .A1(_07640_),
    .A2(_07646_),
    .B1(_05203_),
    .Y(_07648_)
  );
  sg13g2_a21oi_1 _17411_ (
    .A1(addr_i_3_),
    .A2(_00327_),
    .B1(_00605_),
    .Y(_07649_)
  );
  sg13g2_nor2_1 _17412_ (
    .A(_01093_),
    .B(_00559_),
    .Y(_07650_)
  );
  sg13g2_o21ai_1 _17413_ (
    .A1(addr_i_4_),
    .A2(_07649_),
    .B1(_07650_),
    .Y(_07651_)
  );
  sg13g2_a221oi_1 _17414_ (
    .A1(_01758_),
    .A2(_02395_),
    .B1(_07651_),
    .B2(addr_i_5_),
    .C1(_00866_),
    .Y(_07652_)
  );
  sg13g2_nand2_1 _17415_ (
    .A(_00173_),
    .B(_01182_),
    .Y(_07653_)
  );
  sg13g2_a22oi_1 _17416_ (
    .A1(_00408_),
    .A2(_01653_),
    .B1(_00505_),
    .B2(_00491_),
    .Y(_07654_)
  );
  sg13g2_a22oi_1 _17417_ (
    .A1(_09138_),
    .A2(_07653_),
    .B1(_07654_),
    .B2(addr_i_8_),
    .Y(_07655_)
  );
  sg13g2_o21ai_1 _17418_ (
    .A1(addr_i_7_),
    .A2(_07652_),
    .B1(_07655_),
    .Y(_07656_)
  );
  sg13g2_nor2b_1 _17419_ (
    .A(_07648_),
    .B_N(_07656_),
    .Y(_07657_)
  );
  sg13g2_a22oi_1 _17420_ (
    .A1(_01176_),
    .A2(_07637_),
    .B1(_07657_),
    .B2(addr_i_11_),
    .Y(_07659_)
  );
  sg13g2_a221oi_1 _17421_ (
    .A1(addr_i_11_),
    .A2(_07574_),
    .B1(_07616_),
    .B2(_07659_),
    .C1(addr_i_12_),
    .Y(_07660_)
  );
  sg13g2_a21o_1 _17422_ (
    .A1(addr_i_12_),
    .A2(_07490_),
    .B1(_07660_),
    .X(data_o_31_)
  );
  sg13g2_a22oi_1 _17423_ (
    .A1(addr_i_7_),
    .A2(_01815_),
    .B1(_00542_),
    .B2(_01508_),
    .Y(_07661_)
  );
  sg13g2_a21oi_1 _17424_ (
    .A1(_01132_),
    .A2(_01486_),
    .B1(_02368_),
    .Y(_07662_)
  );
  sg13g2_o21ai_1 _17425_ (
    .A1(_00172_),
    .A2(_07661_),
    .B1(_07662_),
    .Y(_07663_)
  );
  sg13g2_a21oi_1 _17426_ (
    .A1(_04063_),
    .A2(_01203_),
    .B1(_00731_),
    .Y(_07664_)
  );
  sg13g2_a21oi_1 _17427_ (
    .A1(_00965_),
    .A2(_00498_),
    .B1(_00020_),
    .Y(_07665_)
  );
  sg13g2_o21ai_1 _17428_ (
    .A1(_07664_),
    .A2(_07665_),
    .B1(addr_i_6_),
    .Y(_07666_)
  );
  sg13g2_o21ai_1 _17429_ (
    .A1(addr_i_7_),
    .A2(_03759_),
    .B1(addr_i_4_),
    .Y(_07667_)
  );
  sg13g2_and2_1 _17430_ (
    .A(_07666_),
    .B(_07667_),
    .X(_07669_)
  );
  sg13g2_nand2b_1 _17431_ (
    .A_N(_04572_),
    .B(_00700_),
    .Y(_07670_)
  );
  sg13g2_nand3_1 _17432_ (
    .A(addr_i_3_),
    .B(_01622_),
    .C(_01222_),
    .Y(_07671_)
  );
  sg13g2_nand3_1 _17433_ (
    .A(_00122_),
    .B(_07670_),
    .C(_07671_),
    .Y(_07672_)
  );
  sg13g2_o21ai_1 _17434_ (
    .A1(_00472_),
    .A2(_09359_),
    .B1(addr_i_7_),
    .Y(_07673_)
  );
  sg13g2_nand3_1 _17435_ (
    .A(addr_i_4_),
    .B(_07672_),
    .C(_07673_),
    .Y(_07674_)
  );
  sg13g2_nor2_1 _17436_ (
    .A(_00473_),
    .B(_00950_),
    .Y(_07675_)
  );
  sg13g2_a21oi_1 _17437_ (
    .A1(_00547_),
    .A2(_00037_),
    .B1(_00020_),
    .Y(_07676_)
  );
  sg13g2_a21oi_1 _17438_ (
    .A1(_04285_),
    .A2(_01004_),
    .B1(_02387_),
    .Y(_07677_)
  );
  sg13g2_or4_1 _17439_ (
    .A(addr_i_4_),
    .B(_07675_),
    .C(_07676_),
    .D(_07677_),
    .X(_07678_)
  );
  sg13g2_a21oi_1 _17440_ (
    .A1(_07674_),
    .A2(_07678_),
    .B1(addr_i_8_),
    .Y(_07680_)
  );
  sg13g2_a22oi_1 _17441_ (
    .A1(addr_i_8_),
    .A2(_07669_),
    .B1(_07680_),
    .B2(addr_i_9_),
    .Y(_07681_)
  );
  sg13g2_a22oi_1 _17442_ (
    .A1(addr_i_9_),
    .A2(_03803_),
    .B1(_07681_),
    .B2(addr_i_10_),
    .Y(_07682_)
  );
  sg13g2_a21oi_1 _17443_ (
    .A1(addr_i_10_),
    .A2(_07663_),
    .B1(_07682_),
    .Y(_07683_)
  );
  sg13g2_o21ai_1 _17444_ (
    .A1(_01103_),
    .A2(_01097_),
    .B1(_07724_),
    .Y(_07684_)
  );
  sg13g2_a22oi_1 _17445_ (
    .A1(addr_i_3_),
    .A2(_06663_),
    .B1(_07684_),
    .B2(addr_i_7_),
    .Y(_07685_)
  );
  sg13g2_nand2_1 _17446_ (
    .A(_02810_),
    .B(_03273_),
    .Y(_07686_)
  );
  sg13g2_a22oi_1 _17447_ (
    .A1(addr_i_6_),
    .A2(_07686_),
    .B1(_02391_),
    .B2(_00779_),
    .Y(_07687_)
  );
  sg13g2_o21ai_1 _17448_ (
    .A1(_07685_),
    .A2(_07687_),
    .B1(addr_i_8_),
    .Y(_07688_)
  );
  sg13g2_nand2_1 _17449_ (
    .A(_00104_),
    .B(_00571_),
    .Y(_07689_)
  );
  sg13g2_a22oi_1 _17450_ (
    .A1(_02404_),
    .A2(_07689_),
    .B1(_00119_),
    .B2(_00778_),
    .Y(_07691_)
  );
  sg13g2_a22oi_1 _17451_ (
    .A1(addr_i_4_),
    .A2(_03662_),
    .B1(_03033_),
    .B2(addr_i_7_),
    .Y(_07692_)
  );
  sg13g2_or3_1 _17452_ (
    .A(_04191_),
    .B(_07691_),
    .C(_07692_),
    .X(_07693_)
  );
  sg13g2_a21oi_1 _17453_ (
    .A1(_02349_),
    .A2(_00317_),
    .B1(_03497_),
    .Y(_07694_)
  );
  sg13g2_a22oi_1 _17454_ (
    .A1(_08399_),
    .A2(_03572_),
    .B1(_07694_),
    .B2(addr_i_8_),
    .Y(_07695_)
  );
  sg13g2_a21oi_1 _17455_ (
    .A1(_07693_),
    .A2(_07695_),
    .B1(addr_i_9_),
    .Y(_07696_)
  );
  sg13g2_nand3_1 _17456_ (
    .A(addr_i_4_),
    .B(_02815_),
    .C(_01060_),
    .Y(_07697_)
  );
  sg13g2_nand2b_1 _17457_ (
    .A_N(_06501_),
    .B(_07697_),
    .Y(_07698_)
  );
  sg13g2_a21oi_1 _17458_ (
    .A1(_00292_),
    .A2(_07698_),
    .B1(addr_i_8_),
    .Y(_07699_)
  );
  sg13g2_nand2_1 _17459_ (
    .A(addr_i_3_),
    .B(_02634_),
    .Y(_07700_)
  );
  sg13g2_nand2_1 _17460_ (
    .A(addr_i_2_),
    .B(_07700_),
    .Y(_07702_)
  );
  sg13g2_a21oi_1 _17461_ (
    .A1(_00443_),
    .A2(_07702_),
    .B1(addr_i_6_),
    .Y(_07703_)
  );
  sg13g2_a21oi_1 _17462_ (
    .A1(_01104_),
    .A2(_03226_),
    .B1(addr_i_3_),
    .Y(_07704_)
  );
  sg13g2_o21ai_1 _17463_ (
    .A1(_07703_),
    .A2(_07704_),
    .B1(addr_i_7_),
    .Y(_07705_)
  );
  sg13g2_nand2_1 _17464_ (
    .A(_06176_),
    .B(_07492_),
    .Y(_07706_)
  );
  sg13g2_a21o_1 _17465_ (
    .A1(_00852_),
    .A2(_01463_),
    .B1(_00445_),
    .X(_07707_)
  );
  sg13g2_nand3_1 _17466_ (
    .A(addr_i_3_),
    .B(addr_i_4_),
    .C(_06473_),
    .Y(_07708_)
  );
  sg13g2_nand3_1 _17467_ (
    .A(_07706_),
    .B(_07707_),
    .C(_07708_),
    .Y(_07709_)
  );
  sg13g2_o21ai_1 _17468_ (
    .A1(_09494_),
    .A2(_02322_),
    .B1(_03288_),
    .Y(_07710_)
  );
  sg13g2_a21oi_1 _17469_ (
    .A1(_03710_),
    .A2(_07710_),
    .B1(_00146_),
    .Y(_07711_)
  );
  sg13g2_o21ai_1 _17470_ (
    .A1(_01380_),
    .A2(_00234_),
    .B1(addr_i_6_),
    .Y(_07714_)
  );
  sg13g2_nand2_1 _17471_ (
    .A(addr_i_8_),
    .B(_07714_),
    .Y(_07715_)
  );
  sg13g2_a22oi_1 _17472_ (
    .A1(addr_i_7_),
    .A2(_07709_),
    .B1(_07711_),
    .B2(_07715_),
    .Y(_07716_)
  );
  sg13g2_a22oi_1 _17473_ (
    .A1(_07699_),
    .A2(_07705_),
    .B1(_00243_),
    .B2(_07716_),
    .Y(_07717_)
  );
  sg13g2_a22oi_1 _17474_ (
    .A1(_07688_),
    .A2(_07696_),
    .B1(_07717_),
    .B2(addr_i_10_),
    .Y(_07718_)
  );
  sg13g2_a21oi_1 _17475_ (
    .A1(_00940_),
    .A2(_04754_),
    .B1(addr_i_5_),
    .Y(_07719_)
  );
  sg13g2_nor2_1 _17476_ (
    .A(_02361_),
    .B(_07719_),
    .Y(_07720_)
  );
  sg13g2_a221oi_1 _17477_ (
    .A1(addr_i_3_),
    .A2(_00827_),
    .B1(_01257_),
    .B2(_01480_),
    .C1(_01794_),
    .Y(_07721_)
  );
  sg13g2_a22oi_1 _17478_ (
    .A1(_01630_),
    .A2(_07720_),
    .B1(_07721_),
    .B2(_02963_),
    .Y(_07722_)
  );
  sg13g2_nor2_1 _17479_ (
    .A(addr_i_7_),
    .B(_07547_),
    .Y(_07723_)
  );
  sg13g2_a21oi_1 _17480_ (
    .A1(_00677_),
    .A2(_03701_),
    .B1(_08011_),
    .Y(_07725_)
  );
  sg13g2_o21ai_1 _17481_ (
    .A1(_02976_),
    .A2(_07001_),
    .B1(_02063_),
    .Y(_07726_)
  );
  sg13g2_o21ai_1 _17482_ (
    .A1(_05603_),
    .A2(_07583_),
    .B1(addr_i_3_),
    .Y(_07727_)
  );
  sg13g2_a21oi_1 _17483_ (
    .A1(_07726_),
    .A2(_07727_),
    .B1(addr_i_6_),
    .Y(_07728_)
  );
  sg13g2_a22oi_1 _17484_ (
    .A1(_03267_),
    .A2(_07723_),
    .B1(_07725_),
    .B2(_07728_),
    .Y(_07729_)
  );
  sg13g2_nor2_1 _17485_ (
    .A(_02368_),
    .B(_07729_),
    .Y(_07730_)
  );
  sg13g2_a22oi_1 _17486_ (
    .A1(_00391_),
    .A2(_03022_),
    .B1(_01611_),
    .B2(_00390_),
    .Y(_07731_)
  );
  sg13g2_o21ai_1 _17487_ (
    .A1(addr_i_2_),
    .A2(_06340_),
    .B1(_01287_),
    .Y(_07732_)
  );
  sg13g2_nand3_1 _17488_ (
    .A(_09487_),
    .B(_02604_),
    .C(_07732_),
    .Y(_07733_)
  );
  sg13g2_nand3b_1 _17489_ (
    .A_N(_07731_),
    .B(_07733_),
    .C(addr_i_10_),
    .Y(_07734_)
  );
  sg13g2_o21ai_1 _17490_ (
    .A1(addr_i_2_),
    .A2(_00011_),
    .B1(addr_i_3_),
    .Y(_07736_)
  );
  sg13g2_a21oi_1 _17491_ (
    .A1(_02528_),
    .A2(_07736_),
    .B1(addr_i_7_),
    .Y(_07737_)
  );
  sg13g2_o21ai_1 _17492_ (
    .A1(_05883_),
    .A2(_07737_),
    .B1(_00084_),
    .Y(_07738_)
  );
  sg13g2_nand2_1 _17493_ (
    .A(addr_i_4_),
    .B(_00702_),
    .Y(_07739_)
  );
  sg13g2_a21oi_1 _17494_ (
    .A1(_00091_),
    .A2(_03089_),
    .B1(_08752_),
    .Y(_07740_)
  );
  sg13g2_a22oi_1 _17495_ (
    .A1(_05062_),
    .A2(_07739_),
    .B1(_07740_),
    .B2(_00351_),
    .Y(_07741_)
  );
  sg13g2_a22oi_1 _17496_ (
    .A1(_06010_),
    .A2(_01551_),
    .B1(_07741_),
    .B2(addr_i_8_),
    .Y(_07742_)
  );
  sg13g2_nor2_1 _17497_ (
    .A(_00226_),
    .B(_05603_),
    .Y(_07743_)
  );
  sg13g2_nand2_1 _17498_ (
    .A(addr_i_4_),
    .B(_06972_),
    .Y(_07744_)
  );
  sg13g2_a22oi_1 _17499_ (
    .A1(addr_i_2_),
    .A2(_07744_),
    .B1(_01127_),
    .B2(addr_i_3_),
    .Y(_07745_)
  );
  sg13g2_a22oi_1 _17500_ (
    .A1(addr_i_3_),
    .A2(_07743_),
    .B1(_07745_),
    .B2(addr_i_6_),
    .Y(_07747_)
  );
  sg13g2_a21o_1 _17501_ (
    .A1(_01453_),
    .A2(_00883_),
    .B1(addr_i_2_),
    .X(_07748_)
  );
  sg13g2_a21oi_1 _17502_ (
    .A1(_02807_),
    .A2(_07748_),
    .B1(_02759_),
    .Y(_07749_)
  );
  sg13g2_a21oi_1 _17503_ (
    .A1(_05517_),
    .A2(_06909_),
    .B1(_00324_),
    .Y(_07750_)
  );
  sg13g2_nor4_1 _17504_ (
    .A(_00113_),
    .B(_07747_),
    .C(_07749_),
    .D(_07750_),
    .Y(_07751_)
  );
  sg13g2_a22oi_1 _17505_ (
    .A1(_07738_),
    .A2(_07742_),
    .B1(_00243_),
    .B2(_07751_),
    .Y(_07752_)
  );
  sg13g2_nor4_1 _17506_ (
    .A(_07722_),
    .B(_07730_),
    .C(_07734_),
    .D(_07752_),
    .Y(_07753_)
  );
  sg13g2_nor2_1 _17507_ (
    .A(_07718_),
    .B(_07753_),
    .Y(_07754_)
  );
  sg13g2_a21oi_1 _17508_ (
    .A1(_04285_),
    .A2(_01738_),
    .B1(_00483_),
    .Y(_07755_)
  );
  sg13g2_o21ai_1 _17509_ (
    .A1(_02935_),
    .A2(_07755_),
    .B1(_01528_),
    .Y(_07756_)
  );
  sg13g2_a21oi_1 _17510_ (
    .A1(_04229_),
    .A2(_07756_),
    .B1(addr_i_6_),
    .Y(_07758_)
  );
  sg13g2_a21oi_1 _17511_ (
    .A1(_00586_),
    .A2(_01462_),
    .B1(_01867_),
    .Y(_07759_)
  );
  sg13g2_a221oi_1 _17512_ (
    .A1(_02976_),
    .A2(_00319_),
    .B1(_01255_),
    .B2(addr_i_7_),
    .C1(_07759_),
    .Y(_07760_)
  );
  sg13g2_nand2_1 _17513_ (
    .A(_00168_),
    .B(_00156_),
    .Y(_07761_)
  );
  sg13g2_o21ai_1 _17514_ (
    .A1(_03263_),
    .A2(_07760_),
    .B1(_07761_),
    .Y(_07762_)
  );
  sg13g2_o21ai_1 _17515_ (
    .A1(_07758_),
    .A2(_07762_),
    .B1(_00367_),
    .Y(_07763_)
  );
  sg13g2_a21oi_1 _17516_ (
    .A1(_00603_),
    .A2(_02533_),
    .B1(_01114_),
    .Y(_07764_)
  );
  sg13g2_a22oi_1 _17517_ (
    .A1(_02277_),
    .A2(_07157_),
    .B1(_07764_),
    .B2(_03526_),
    .Y(_07765_)
  );
  sg13g2_a21oi_1 _17518_ (
    .A1(_00370_),
    .A2(_01625_),
    .B1(addr_i_2_),
    .Y(_07766_)
  );
  sg13g2_a21o_1 _17519_ (
    .A1(addr_i_4_),
    .A2(_03932_),
    .B1(_07766_),
    .X(_07767_)
  );
  sg13g2_nor2_1 _17520_ (
    .A(_00676_),
    .B(_06541_),
    .Y(_07769_)
  );
  sg13g2_a21oi_1 _17521_ (
    .A1(_07769_),
    .A2(_04371_),
    .B1(addr_i_3_),
    .Y(_07770_)
  );
  sg13g2_a221oi_1 _17522_ (
    .A1(_08388_),
    .A2(_00282_),
    .B1(_07767_),
    .B2(addr_i_3_),
    .C1(_07770_),
    .Y(_07771_)
  );
  sg13g2_nor2_1 _17523_ (
    .A(_08674_),
    .B(_07771_),
    .Y(_07772_)
  );
  sg13g2_nor3_1 _17524_ (
    .A(addr_i_9_),
    .B(_07765_),
    .C(_07772_),
    .Y(_07773_)
  );
  sg13g2_nor2_1 _17525_ (
    .A(_02777_),
    .B(_00227_),
    .Y(_07774_)
  );
  sg13g2_nor3_1 _17526_ (
    .A(addr_i_6_),
    .B(_03308_),
    .C(_04939_),
    .Y(_07775_)
  );
  sg13g2_a22oi_1 _17527_ (
    .A1(_00816_),
    .A2(_07774_),
    .B1(_07775_),
    .B2(_00860_),
    .Y(_07776_)
  );
  sg13g2_a22oi_1 _17528_ (
    .A1(addr_i_4_),
    .A2(_02585_),
    .B1(_06264_),
    .B2(addr_i_3_),
    .Y(_07777_)
  );
  sg13g2_a21oi_1 _17529_ (
    .A1(_00155_),
    .A2(_07458_),
    .B1(_07777_),
    .Y(_07778_)
  );
  sg13g2_a21oi_1 _17530_ (
    .A1(_09260_),
    .A2(_02032_),
    .B1(addr_i_4_),
    .Y(_07780_)
  );
  sg13g2_nor3_1 _17531_ (
    .A(_07514_),
    .B(_07778_),
    .C(_07780_),
    .Y(_07781_)
  );
  sg13g2_nand2_1 _17532_ (
    .A(addr_i_3_),
    .B(_07025_),
    .Y(_07782_)
  );
  sg13g2_a21oi_1 _17533_ (
    .A1(_00739_),
    .A2(_07782_),
    .B1(addr_i_4_),
    .Y(_07783_)
  );
  sg13g2_a221oi_1 _17534_ (
    .A1(_00838_),
    .A2(_03556_),
    .B1(_03401_),
    .B2(_00999_),
    .C1(_07783_),
    .Y(_07784_)
  );
  sg13g2_nor2_1 _17535_ (
    .A(_01099_),
    .B(_07784_),
    .Y(_07785_)
  );
  sg13g2_o21ai_1 _17536_ (
    .A1(_01277_),
    .A2(_01815_),
    .B1(_07934_),
    .Y(_07786_)
  );
  sg13g2_nand3_1 _17537_ (
    .A(_00749_),
    .B(_00771_),
    .C(_01912_),
    .Y(_07787_)
  );
  sg13g2_o21ai_1 _17538_ (
    .A1(_07786_),
    .A2(_07787_),
    .B1(addr_i_9_),
    .Y(_07788_)
  );
  sg13g2_nor4_1 _17539_ (
    .A(_07776_),
    .B(_07781_),
    .C(_07785_),
    .D(_07788_),
    .Y(_07789_)
  );
  sg13g2_a22oi_1 _17540_ (
    .A1(_07763_),
    .A2(_07773_),
    .B1(_07789_),
    .B2(_01773_),
    .Y(_07791_)
  );
  sg13g2_nor3_1 _17541_ (
    .A(_00715_),
    .B(_00491_),
    .C(_01216_),
    .Y(_07792_)
  );
  sg13g2_o21ai_1 _17542_ (
    .A1(addr_i_2_),
    .A2(_02514_),
    .B1(_01114_),
    .Y(_07793_)
  );
  sg13g2_a21oi_1 _17543_ (
    .A1(_01104_),
    .A2(_07793_),
    .B1(_03132_),
    .Y(_07794_)
  );
  sg13g2_a22oi_1 _17544_ (
    .A1(_04969_),
    .A2(_07792_),
    .B1(_07794_),
    .B2(_02700_),
    .Y(_07795_)
  );
  sg13g2_nor2_1 _17545_ (
    .A(_08166_),
    .B(_00280_),
    .Y(_07796_)
  );
  sg13g2_o21ai_1 _17546_ (
    .A1(addr_i_3_),
    .A2(_00574_),
    .B1(_07796_),
    .Y(_07797_)
  );
  sg13g2_a21oi_1 _17547_ (
    .A1(_07768_),
    .A2(_01037_),
    .B1(addr_i_2_),
    .Y(_07798_)
  );
  sg13g2_a22oi_1 _17548_ (
    .A1(addr_i_2_),
    .A2(_07797_),
    .B1(_07798_),
    .B2(_07554_),
    .Y(_07799_)
  );
  sg13g2_nor2_1 _17549_ (
    .A(_08674_),
    .B(_07799_),
    .Y(_07800_)
  );
  sg13g2_nor2_1 _17550_ (
    .A(_08464_),
    .B(_02184_),
    .Y(_07802_)
  );
  sg13g2_a21oi_1 _17551_ (
    .A1(_00227_),
    .A2(_00333_),
    .B1(_07802_),
    .Y(_07803_)
  );
  sg13g2_a21o_1 _17552_ (
    .A1(_02250_),
    .A2(_04186_),
    .B1(_05281_),
    .X(_07804_)
  );
  sg13g2_a21oi_1 _17553_ (
    .A1(_00545_),
    .A2(_07804_),
    .B1(_04041_),
    .Y(_07805_)
  );
  sg13g2_a22oi_1 _17554_ (
    .A1(_01881_),
    .A2(_03045_),
    .B1(_07805_),
    .B2(addr_i_7_),
    .Y(_07806_)
  );
  sg13g2_a22oi_1 _17555_ (
    .A1(addr_i_7_),
    .A2(_07803_),
    .B1(_07806_),
    .B2(addr_i_8_),
    .Y(_07807_)
  );
  sg13g2_nor2_1 _17556_ (
    .A(_07800_),
    .B(_07807_),
    .Y(_07808_)
  );
  sg13g2_a21oi_1 _17557_ (
    .A1(_00383_),
    .A2(_00242_),
    .B1(_03523_),
    .Y(_07809_)
  );
  sg13g2_o21ai_1 _17558_ (
    .A1(addr_i_3_),
    .A2(_07809_),
    .B1(_00655_),
    .Y(_07810_)
  );
  sg13g2_nor3_1 _17559_ (
    .A(addr_i_6_),
    .B(_04307_),
    .C(_00099_),
    .Y(_07811_)
  );
  sg13g2_o21ai_1 _17560_ (
    .A1(_05575_),
    .A2(_07811_),
    .B1(addr_i_5_),
    .Y(_07813_)
  );
  sg13g2_nand3_1 _17561_ (
    .A(_06143_),
    .B(_00086_),
    .C(_08520_),
    .Y(_07814_)
  );
  sg13g2_a21oi_1 _17562_ (
    .A1(_07813_),
    .A2(_07814_),
    .B1(_09491_),
    .Y(_07815_)
  );
  sg13g2_o21ai_1 _17563_ (
    .A1(addr_i_4_),
    .A2(_00242_),
    .B1(_08741_),
    .Y(_07816_)
  );
  sg13g2_a22oi_1 _17564_ (
    .A1(_00381_),
    .A2(_07816_),
    .B1(addr_i_2_),
    .B2(addr_i_7_),
    .Y(_07817_)
  );
  sg13g2_a22oi_1 _17565_ (
    .A1(addr_i_2_),
    .A2(_07810_),
    .B1(_07815_),
    .B2(_07817_),
    .Y(_07818_)
  );
  sg13g2_nor2_1 _17566_ (
    .A(_06695_),
    .B(_07818_),
    .Y(_07819_)
  );
  sg13g2_a21oi_1 _17567_ (
    .A1(_02077_),
    .A2(_01841_),
    .B1(_04041_),
    .Y(_07820_)
  );
  sg13g2_a21oi_1 _17568_ (
    .A1(_00671_),
    .A2(_02187_),
    .B1(addr_i_3_),
    .Y(_07821_)
  );
  sg13g2_a22oi_1 _17569_ (
    .A1(_00594_),
    .A2(_02203_),
    .B1(_07820_),
    .B2(_07821_),
    .Y(_07822_)
  );
  sg13g2_nand2b_1 _17570_ (
    .A_N(_01735_),
    .B(_05979_),
    .Y(_07825_)
  );
  sg13g2_a221oi_1 _17571_ (
    .A1(_08056_),
    .A2(_02289_),
    .B1(_07825_),
    .B2(addr_i_6_),
    .C1(addr_i_7_),
    .Y(_07826_)
  );
  sg13g2_a22oi_1 _17572_ (
    .A1(addr_i_7_),
    .A2(_07822_),
    .B1(_07826_),
    .B2(addr_i_8_),
    .Y(_07827_)
  );
  sg13g2_nor3_1 _17573_ (
    .A(addr_i_9_),
    .B(_07819_),
    .C(_07827_),
    .Y(_07828_)
  );
  sg13g2_a22oi_1 _17574_ (
    .A1(_07795_),
    .A2(_07808_),
    .B1(addr_i_10_),
    .B2(_07828_),
    .Y(_07829_)
  );
  sg13g2_or2_1 _17575_ (
    .A(_07791_),
    .B(_07829_),
    .X(_07830_)
  );
  sg13g2_a21oi_1 _17576_ (
    .A1(addr_i_2_),
    .A2(_00418_),
    .B1(_00713_),
    .Y(_07831_)
  );
  sg13g2_o21ai_1 _17577_ (
    .A1(_00648_),
    .A2(_07831_),
    .B1(_06206_),
    .Y(_07832_)
  );
  sg13g2_nor3_1 _17578_ (
    .A(addr_i_5_),
    .B(_05490_),
    .C(_07603_),
    .Y(_07833_)
  );
  sg13g2_a21o_1 _17579_ (
    .A1(_01571_),
    .A2(_07832_),
    .B1(_07833_),
    .X(_07834_)
  );
  sg13g2_a21oi_1 _17580_ (
    .A1(_00287_),
    .A2(_05263_),
    .B1(_00032_),
    .Y(_07836_)
  );
  sg13g2_a21oi_1 _17581_ (
    .A1(_05501_),
    .A2(_00301_),
    .B1(_07836_),
    .Y(_07837_)
  );
  sg13g2_o21ai_1 _17582_ (
    .A1(addr_i_8_),
    .A2(_07837_),
    .B1(addr_i_9_),
    .Y(_07838_)
  );
  sg13g2_o21ai_1 _17583_ (
    .A1(_03523_),
    .A2(_01869_),
    .B1(addr_i_2_),
    .Y(_07839_)
  );
  sg13g2_a22oi_1 _17584_ (
    .A1(_05427_),
    .A2(_07839_),
    .B1(addr_i_3_),
    .B2(_07403_),
    .Y(_07840_)
  );
  sg13g2_a22oi_1 _17585_ (
    .A1(_02257_),
    .A2(_07834_),
    .B1(_07838_),
    .B2(_07840_),
    .Y(_07841_)
  );
  sg13g2_a22oi_1 _17586_ (
    .A1(addr_i_4_),
    .A2(_03045_),
    .B1(_06519_),
    .B2(addr_i_8_),
    .Y(_07842_)
  );
  sg13g2_a22oi_1 _17587_ (
    .A1(_02173_),
    .A2(_00960_),
    .B1(_04679_),
    .B2(_06684_),
    .Y(_07843_)
  );
  sg13g2_nor3_1 _17588_ (
    .A(_01517_),
    .B(_07842_),
    .C(_07843_),
    .Y(_07844_)
  );
  sg13g2_nand2_1 _17589_ (
    .A(addr_i_3_),
    .B(_02525_),
    .Y(_07845_)
  );
  sg13g2_a21oi_1 _17590_ (
    .A1(_07569_),
    .A2(_07845_),
    .B1(addr_i_5_),
    .Y(_07847_)
  );
  sg13g2_nor2_1 _17591_ (
    .A(_01746_),
    .B(_07847_),
    .Y(_07848_)
  );
  sg13g2_nor2_1 _17592_ (
    .A(_07945_),
    .B(_07848_),
    .Y(_07849_)
  );
  sg13g2_nand3_1 _17593_ (
    .A(addr_i_2_),
    .B(_02383_),
    .C(_00785_),
    .Y(_07850_)
  );
  sg13g2_nand3_1 _17594_ (
    .A(_03919_),
    .B(_00371_),
    .C(_04765_),
    .Y(_07851_)
  );
  sg13g2_nand3_1 _17595_ (
    .A(_05218_),
    .B(_07850_),
    .C(_07851_),
    .Y(_07852_)
  );
  sg13g2_nand2_1 _17596_ (
    .A(_09507_),
    .B(_00499_),
    .Y(_07853_)
  );
  sg13g2_a21oi_1 _17597_ (
    .A1(_07852_),
    .A2(_07853_),
    .B1(addr_i_8_),
    .Y(_07854_)
  );
  sg13g2_nor4_1 _17598_ (
    .A(addr_i_9_),
    .B(_07844_),
    .C(_07849_),
    .D(_07854_),
    .Y(_07855_)
  );
  sg13g2_o21ai_1 _17599_ (
    .A1(_07841_),
    .A2(_07855_),
    .B1(addr_i_10_),
    .Y(_07856_)
  );
  sg13g2_a21oi_1 _17600_ (
    .A1(addr_i_2_),
    .A2(_00786_),
    .B1(_01779_),
    .Y(_07858_)
  );
  sg13g2_o21ai_1 _17601_ (
    .A1(addr_i_3_),
    .A2(_07858_),
    .B1(_03581_),
    .Y(_07859_)
  );
  sg13g2_nand2_1 _17602_ (
    .A(_00827_),
    .B(_01309_),
    .Y(_07860_)
  );
  sg13g2_o21ai_1 _17603_ (
    .A1(_05557_),
    .A2(_01309_),
    .B1(_07860_),
    .Y(_07861_)
  );
  sg13g2_a22oi_1 _17604_ (
    .A1(addr_i_2_),
    .A2(_00498_),
    .B1(_03348_),
    .B2(_02569_),
    .Y(_07862_)
  );
  sg13g2_or2_1 _17605_ (
    .A(addr_i_8_),
    .B(_07862_),
    .X(_07863_)
  );
  sg13g2_a221oi_1 _17606_ (
    .A1(addr_i_7_),
    .A2(_07859_),
    .B1(_07861_),
    .B2(_00402_),
    .C1(_07863_),
    .Y(_07864_)
  );
  sg13g2_nor2_1 _17607_ (
    .A(_00032_),
    .B(_04261_),
    .Y(_07865_)
  );
  sg13g2_nand2b_1 _17608_ (
    .A_N(_06179_),
    .B(_07865_),
    .Y(_07866_)
  );
  sg13g2_nand3_1 _17609_ (
    .A(_00428_),
    .B(_01007_),
    .C(_00712_),
    .Y(_07867_)
  );
  sg13g2_nand3_1 _17610_ (
    .A(addr_i_8_),
    .B(_07866_),
    .C(_07867_),
    .Y(_07869_)
  );
  sg13g2_o21ai_1 _17611_ (
    .A1(addr_i_3_),
    .A2(_00591_),
    .B1(_00778_),
    .Y(_07870_)
  );
  sg13g2_a21oi_1 _17612_ (
    .A1(addr_i_4_),
    .A2(addr_i_6_),
    .B1(addr_i_2_),
    .Y(_07871_)
  );
  sg13g2_nand2_1 _17613_ (
    .A(_00046_),
    .B(_07871_),
    .Y(_07872_)
  );
  sg13g2_a21oi_1 _17614_ (
    .A1(_00603_),
    .A2(_07872_),
    .B1(addr_i_5_),
    .Y(_07873_)
  );
  sg13g2_nor3_1 _17615_ (
    .A(_04613_),
    .B(_07870_),
    .C(_07873_),
    .Y(_07874_)
  );
  sg13g2_o21ai_1 _17616_ (
    .A1(_07869_),
    .A2(_07874_),
    .B1(addr_i_9_),
    .Y(_07875_)
  );
  sg13g2_nand2_1 _17617_ (
    .A(_00157_),
    .B(_07025_),
    .Y(_07876_)
  );
  sg13g2_o21ai_1 _17618_ (
    .A1(_01292_),
    .A2(_04837_),
    .B1(addr_i_3_),
    .Y(_07877_)
  );
  sg13g2_o21ai_1 _17619_ (
    .A1(_01837_),
    .A2(_00279_),
    .B1(addr_i_4_),
    .Y(_07878_)
  );
  sg13g2_nand3_1 _17620_ (
    .A(_07876_),
    .B(_07877_),
    .C(_07878_),
    .Y(_07880_)
  );
  sg13g2_nor3_1 _17621_ (
    .A(_01970_),
    .B(_00343_),
    .C(_00840_),
    .Y(_07881_)
  );
  sg13g2_nor2_1 _17622_ (
    .A(_01746_),
    .B(_07881_),
    .Y(_07882_)
  );
  sg13g2_nor3_1 _17623_ (
    .A(_01481_),
    .B(_01611_),
    .C(_07882_),
    .Y(_07883_)
  );
  sg13g2_a22oi_1 _17624_ (
    .A1(_03374_),
    .A2(_07880_),
    .B1(_07883_),
    .B2(addr_i_10_),
    .Y(_07884_)
  );
  sg13g2_o21ai_1 _17625_ (
    .A1(_07864_),
    .A2(_07875_),
    .B1(_07884_),
    .Y(_07885_)
  );
  sg13g2_and2_1 _17626_ (
    .A(_07856_),
    .B(_07885_),
    .X(_07886_)
  );
  sg13g2_mux4_1 _17627_ (
    .A0(_07683_),
    .A1(_07754_),
    .A2(_07830_),
    .A3(_07886_),
    .S0(_03051_),
    .S1(_02251_),
    .X(data_o_3_)
  );
  sg13g2_nand2_1 _17628_ (
    .A(_00138_),
    .B(_01432_),
    .Y(_07887_)
  );
  sg13g2_a21oi_1 _17629_ (
    .A1(_00482_),
    .A2(_00702_),
    .B1(_09513_),
    .Y(_07888_)
  );
  sg13g2_a22oi_1 _17630_ (
    .A1(_00258_),
    .A2(_07887_),
    .B1(_07888_),
    .B2(_02026_),
    .Y(_07890_)
  );
  sg13g2_o21ai_1 _17631_ (
    .A1(_02744_),
    .A2(_03485_),
    .B1(_07890_),
    .Y(_07891_)
  );
  sg13g2_a21oi_1 _17632_ (
    .A1(_01453_),
    .A2(_07700_),
    .B1(_02012_),
    .Y(_07892_)
  );
  sg13g2_a22oi_1 _17633_ (
    .A1(_01019_),
    .A2(_06276_),
    .B1(_04837_),
    .B2(_07892_),
    .Y(_07893_)
  );
  sg13g2_o21ai_1 _17634_ (
    .A1(_07614_),
    .A2(_07893_),
    .B1(addr_i_9_),
    .Y(_07894_)
  );
  sg13g2_a21oi_1 _17635_ (
    .A1(_05435_),
    .A2(_04195_),
    .B1(addr_i_4_),
    .Y(_07895_)
  );
  sg13g2_o21ai_1 _17636_ (
    .A1(_09513_),
    .A2(_02626_),
    .B1(_03519_),
    .Y(_07896_)
  );
  sg13g2_nor4_1 _17637_ (
    .A(_01281_),
    .B(_01986_),
    .C(_07895_),
    .D(_07896_),
    .Y(_07897_)
  );
  sg13g2_nor2_1 _17638_ (
    .A(_09205_),
    .B(_01097_),
    .Y(_07898_)
  );
  sg13g2_a21oi_1 _17639_ (
    .A1(_01473_),
    .A2(_00567_),
    .B1(addr_i_3_),
    .Y(_07899_)
  );
  sg13g2_o21ai_1 _17640_ (
    .A1(_07898_),
    .A2(_07899_),
    .B1(_00276_),
    .Y(_07901_)
  );
  sg13g2_o21ai_1 _17641_ (
    .A1(_08487_),
    .A2(_07897_),
    .B1(_07901_),
    .Y(_07902_)
  );
  sg13g2_a22oi_1 _17642_ (
    .A1(_01119_),
    .A2(_07891_),
    .B1(_07894_),
    .B2(_07902_),
    .Y(_07903_)
  );
  sg13g2_nor3_1 _17643_ (
    .A(_01472_),
    .B(_07658_),
    .C(_00961_),
    .Y(_07904_)
  );
  sg13g2_nor2_1 _17644_ (
    .A(_01016_),
    .B(_07904_),
    .Y(_07905_)
  );
  sg13g2_nor3_1 _17645_ (
    .A(_00096_),
    .B(_04400_),
    .C(_04316_),
    .Y(_07906_)
  );
  sg13g2_a21oi_1 _17646_ (
    .A1(_07905_),
    .A2(_07906_),
    .B1(_00949_),
    .Y(_07907_)
  );
  sg13g2_a21oi_1 _17647_ (
    .A1(_00441_),
    .A2(_02136_),
    .B1(addr_i_3_),
    .Y(_07908_)
  );
  sg13g2_o21ai_1 _17648_ (
    .A1(_09094_),
    .A2(_07908_),
    .B1(_06717_),
    .Y(_07909_)
  );
  sg13g2_o21ai_1 _17649_ (
    .A1(_03993_),
    .A2(_03648_),
    .B1(_09499_),
    .Y(_07910_)
  );
  sg13g2_nand3b_1 _17650_ (
    .A_N(_07907_),
    .B(_07909_),
    .C(_07910_),
    .Y(_07912_)
  );
  sg13g2_o21ai_1 _17651_ (
    .A1(_08343_),
    .A2(_06950_),
    .B1(addr_i_3_),
    .Y(_07913_)
  );
  sg13g2_nand3_1 _17652_ (
    .A(_09491_),
    .B(addr_i_4_),
    .C(_01738_),
    .Y(_07914_)
  );
  sg13g2_nand4_1 _17653_ (
    .A(_00476_),
    .B(_00250_),
    .C(_07913_),
    .D(_07914_),
    .Y(_07915_)
  );
  sg13g2_a22oi_1 _17654_ (
    .A1(_00861_),
    .A2(_00574_),
    .B1(_03980_),
    .B2(_03033_),
    .Y(_07916_)
  );
  sg13g2_o21ai_1 _17655_ (
    .A1(addr_i_7_),
    .A2(_00692_),
    .B1(_01570_),
    .Y(_07917_)
  );
  sg13g2_a22oi_1 _17656_ (
    .A1(addr_i_4_),
    .A2(_07917_),
    .B1(_03455_),
    .B2(addr_i_8_),
    .Y(_07918_)
  );
  sg13g2_o21ai_1 _17657_ (
    .A1(_01615_),
    .A2(_07916_),
    .B1(_07918_),
    .Y(_07919_)
  );
  sg13g2_a21oi_1 _17658_ (
    .A1(addr_i_6_),
    .A2(_07915_),
    .B1(_07919_),
    .Y(_07920_)
  );
  sg13g2_a22oi_1 _17659_ (
    .A1(addr_i_8_),
    .A2(_07912_),
    .B1(_07920_),
    .B2(addr_i_9_),
    .Y(_07921_)
  );
  sg13g2_nor2_1 _17660_ (
    .A(_07903_),
    .B(_07921_),
    .Y(_07923_)
  );
  sg13g2_o21ai_1 _17661_ (
    .A1(_05711_),
    .A2(_00901_),
    .B1(_00020_),
    .Y(_07924_)
  );
  sg13g2_nor3_1 _17662_ (
    .A(_00927_),
    .B(_07812_),
    .C(_00158_),
    .Y(_07925_)
  );
  sg13g2_a22oi_1 _17663_ (
    .A1(addr_i_7_),
    .A2(_07924_),
    .B1(_07925_),
    .B2(_02361_),
    .Y(_07926_)
  );
  sg13g2_nand2_1 _17664_ (
    .A(_01384_),
    .B(_00998_),
    .Y(_07927_)
  );
  sg13g2_nand3_1 _17665_ (
    .A(_07779_),
    .B(_01432_),
    .C(_07927_),
    .Y(_07928_)
  );
  sg13g2_a221oi_1 _17666_ (
    .A1(_00666_),
    .A2(_00645_),
    .B1(_07928_),
    .B2(_04068_),
    .C1(_09271_),
    .Y(_07929_)
  );
  sg13g2_a21oi_1 _17667_ (
    .A1(_08399_),
    .A2(_07926_),
    .B1(_07929_),
    .Y(_07930_)
  );
  sg13g2_a21oi_1 _17668_ (
    .A1(_04162_),
    .A2(_02799_),
    .B1(addr_i_6_),
    .Y(_07931_)
  );
  sg13g2_o21ai_1 _17669_ (
    .A1(_08896_),
    .A2(_03172_),
    .B1(addr_i_4_),
    .Y(_07932_)
  );
  sg13g2_a21oi_1 _17670_ (
    .A1(_00671_),
    .A2(_07932_),
    .B1(addr_i_7_),
    .Y(_07935_)
  );
  sg13g2_o21ai_1 _17671_ (
    .A1(_07931_),
    .A2(_07935_),
    .B1(_02271_),
    .Y(_07936_)
  );
  sg13g2_a21oi_1 _17672_ (
    .A1(_06032_),
    .A2(_00358_),
    .B1(addr_i_5_),
    .Y(_07937_)
  );
  sg13g2_a21oi_1 _17673_ (
    .A1(_00716_),
    .A2(_00907_),
    .B1(_02990_),
    .Y(_07938_)
  );
  sg13g2_o21ai_1 _17674_ (
    .A1(_07937_),
    .A2(_07938_),
    .B1(addr_i_7_),
    .Y(_07939_)
  );
  sg13g2_nand4_1 _17675_ (
    .A(_01043_),
    .B(_02052_),
    .C(_07936_),
    .D(_07939_),
    .Y(_07940_)
  );
  sg13g2_o21ai_1 _17676_ (
    .A1(_07293_),
    .A2(_07930_),
    .B1(_07940_),
    .Y(_07941_)
  );
  sg13g2_a21oi_1 _17677_ (
    .A1(addr_i_7_),
    .A2(_07480_),
    .B1(_02154_),
    .Y(_07942_)
  );
  sg13g2_nand2_1 _17678_ (
    .A(_03314_),
    .B(_02283_),
    .Y(_07943_)
  );
  sg13g2_a21oi_1 _17679_ (
    .A1(addr_i_2_),
    .A2(_07943_),
    .B1(_03643_),
    .Y(_07944_)
  );
  sg13g2_o21ai_1 _17680_ (
    .A1(addr_i_4_),
    .A2(_07942_),
    .B1(_07944_),
    .Y(_07946_)
  );
  sg13g2_a21oi_1 _17681_ (
    .A1(_00435_),
    .A2(_00413_),
    .B1(addr_i_4_),
    .Y(_07947_)
  );
  sg13g2_o21ai_1 _17682_ (
    .A1(_00209_),
    .A2(_07947_),
    .B1(addr_i_3_),
    .Y(_07948_)
  );
  sg13g2_nand2_1 _17683_ (
    .A(addr_i_8_),
    .B(_07948_),
    .Y(_07949_)
  );
  sg13g2_nor3_1 _17684_ (
    .A(_02330_),
    .B(_02361_),
    .C(_04316_),
    .Y(_07950_)
  );
  sg13g2_nor2_1 _17685_ (
    .A(_04384_),
    .B(_08453_),
    .Y(_07951_)
  );
  sg13g2_nor4_1 _17686_ (
    .A(_01127_),
    .B(_07951_),
    .C(_03149_),
    .D(_07054_),
    .Y(_07952_)
  );
  sg13g2_a21oi_1 _17687_ (
    .A1(_07950_),
    .A2(_07952_),
    .B1(_00659_),
    .Y(_07953_)
  );
  sg13g2_a22oi_1 _17688_ (
    .A1(_00116_),
    .A2(_07946_),
    .B1(_07949_),
    .B2(_07953_),
    .Y(_07954_)
  );
  sg13g2_nand3_1 _17689_ (
    .A(_05648_),
    .B(_00739_),
    .C(_04943_),
    .Y(_07955_)
  );
  sg13g2_a21oi_1 _17690_ (
    .A1(_05391_),
    .A2(_01230_),
    .B1(addr_i_4_),
    .Y(_07957_)
  );
  sg13g2_a22oi_1 _17691_ (
    .A1(addr_i_4_),
    .A2(_07955_),
    .B1(_07957_),
    .B2(_02361_),
    .Y(_07958_)
  );
  sg13g2_nor2_1 _17692_ (
    .A(_00802_),
    .B(_07958_),
    .Y(_07959_)
  );
  sg13g2_nand3_1 _17693_ (
    .A(addr_i_6_),
    .B(_03954_),
    .C(_03371_),
    .Y(_07960_)
  );
  sg13g2_o21ai_1 _17694_ (
    .A1(_03648_),
    .A2(_00797_),
    .B1(_07960_),
    .Y(_07961_)
  );
  sg13g2_o21ai_1 _17695_ (
    .A1(_07614_),
    .A2(_07961_),
    .B1(addr_i_9_),
    .Y(_07962_)
  );
  sg13g2_nor3_1 _17696_ (
    .A(_07954_),
    .B(_07959_),
    .C(_07962_),
    .Y(_07963_)
  );
  sg13g2_a22oi_1 _17697_ (
    .A1(_09326_),
    .A2(_07941_),
    .B1(_07963_),
    .B2(_03841_),
    .Y(_07964_)
  );
  sg13g2_a22oi_1 _17698_ (
    .A1(_01774_),
    .A2(_07923_),
    .B1(_07964_),
    .B2(addr_i_11_),
    .Y(_07965_)
  );
  sg13g2_a21oi_1 _17699_ (
    .A1(_06784_),
    .A2(_00405_),
    .B1(_01114_),
    .Y(_07966_)
  );
  sg13g2_o21ai_1 _17700_ (
    .A1(_05603_),
    .A2(_07966_),
    .B1(_08011_),
    .Y(_07968_)
  );
  sg13g2_nand2_1 _17701_ (
    .A(_00785_),
    .B(_01967_),
    .Y(_07969_)
  );
  sg13g2_a22oi_1 _17702_ (
    .A1(addr_i_2_),
    .A2(_07969_),
    .B1(_01567_),
    .B2(addr_i_3_),
    .Y(_07970_)
  );
  sg13g2_nor3_1 _17703_ (
    .A(addr_i_7_),
    .B(_01459_),
    .C(_00743_),
    .Y(_07971_)
  );
  sg13g2_a21oi_1 _17704_ (
    .A1(_00482_),
    .A2(_00618_),
    .B1(_00083_),
    .Y(_07972_)
  );
  sg13g2_a22oi_1 _17705_ (
    .A1(_02803_),
    .A2(_07971_),
    .B1(_07972_),
    .B2(_01935_),
    .Y(_07973_)
  );
  sg13g2_a21oi_1 _17706_ (
    .A1(_07968_),
    .A2(_07970_),
    .B1(_07973_),
    .Y(_07974_)
  );
  sg13g2_nor3_1 _17707_ (
    .A(addr_i_8_),
    .B(_07171_),
    .C(_07974_),
    .Y(_07975_)
  );
  sg13g2_a21oi_1 _17708_ (
    .A1(_00688_),
    .A2(_07288_),
    .B1(_00067_),
    .Y(_07976_)
  );
  sg13g2_a21oi_1 _17709_ (
    .A1(_01103_),
    .A2(_04943_),
    .B1(addr_i_4_),
    .Y(_07977_)
  );
  sg13g2_nor3_1 _17710_ (
    .A(addr_i_3_),
    .B(_09271_),
    .C(_00022_),
    .Y(_07979_)
  );
  sg13g2_nor2_1 _17711_ (
    .A(_07558_),
    .B(_01765_),
    .Y(_07980_)
  );
  sg13g2_nor4_1 _17712_ (
    .A(_07976_),
    .B(_07977_),
    .C(_07979_),
    .D(_07980_),
    .Y(_07981_)
  );
  sg13g2_o21ai_1 _17713_ (
    .A1(_01391_),
    .A2(_07981_),
    .B1(_01374_),
    .Y(_07982_)
  );
  sg13g2_nor2_1 _17714_ (
    .A(_04152_),
    .B(_01360_),
    .Y(_07983_)
  );
  sg13g2_a21oi_1 _17715_ (
    .A1(addr_i_9_),
    .A2(_07983_),
    .B1(addr_i_10_),
    .Y(_07984_)
  );
  sg13g2_o21ai_1 _17716_ (
    .A1(_07975_),
    .A2(_07982_),
    .B1(_07984_),
    .Y(_07985_)
  );
  sg13g2_nand2_1 _17717_ (
    .A(addr_i_7_),
    .B(_03745_),
    .Y(_07986_)
  );
  sg13g2_nor2_1 _17718_ (
    .A(_00807_),
    .B(_01357_),
    .Y(_07987_)
  );
  sg13g2_o21ai_1 _17719_ (
    .A1(_05974_),
    .A2(_07986_),
    .B1(_07987_),
    .Y(_07988_)
  );
  sg13g2_nand3_1 _17720_ (
    .A(addr_i_11_),
    .B(_07985_),
    .C(_07988_),
    .Y(_07990_)
  );
  sg13g2_nand2b_1 _17721_ (
    .A_N(_07965_),
    .B(_07990_),
    .Y(_07991_)
  );
  sg13g2_nor2_1 _17722_ (
    .A(_00100_),
    .B(_00087_),
    .Y(_07992_)
  );
  sg13g2_a21oi_1 _17723_ (
    .A1(_00103_),
    .A2(_00007_),
    .B1(addr_i_4_),
    .Y(_07993_)
  );
  sg13g2_a21oi_1 _17724_ (
    .A1(addr_i_4_),
    .A2(_07992_),
    .B1(_07993_),
    .Y(_07994_)
  );
  sg13g2_nand3_1 _17725_ (
    .A(addr_i_4_),
    .B(_04396_),
    .C(_01257_),
    .Y(_07995_)
  );
  sg13g2_a21oi_1 _17726_ (
    .A1(_03420_),
    .A2(_07995_),
    .B1(_01279_),
    .Y(_07996_)
  );
  sg13g2_a21oi_1 _17727_ (
    .A1(_01324_),
    .A2(_07994_),
    .B1(_07996_),
    .Y(_07997_)
  );
  sg13g2_nor2_1 _17728_ (
    .A(addr_i_5_),
    .B(_09501_),
    .Y(_07998_)
  );
  sg13g2_a22oi_1 _17729_ (
    .A1(_00183_),
    .A2(_00414_),
    .B1(_01754_),
    .B2(_01320_),
    .Y(_07999_)
  );
  sg13g2_nor2_1 _17730_ (
    .A(_01279_),
    .B(_07999_),
    .Y(_08001_)
  );
  sg13g2_a22oi_1 _17731_ (
    .A1(_02268_),
    .A2(_07998_),
    .B1(_08001_),
    .B2(_00061_),
    .Y(_08002_)
  );
  sg13g2_a22oi_1 _17732_ (
    .A1(_00048_),
    .A2(_07997_),
    .B1(_08002_),
    .B2(_01612_),
    .Y(_08003_)
  );
  sg13g2_inv_1 _17733_ (
    .A(_08003_),
    .Y(_08004_)
  );
  sg13g2_a22oi_1 _17734_ (
    .A1(addr_i_4_),
    .A2(_00808_),
    .B1(_01825_),
    .B2(_07215_),
    .Y(_08005_)
  );
  sg13g2_o21ai_1 _17735_ (
    .A1(_06740_),
    .A2(_01127_),
    .B1(_06806_),
    .Y(_08006_)
  );
  sg13g2_o21ai_1 _17736_ (
    .A1(addr_i_5_),
    .A2(_08005_),
    .B1(_08006_),
    .Y(_08007_)
  );
  sg13g2_and2_1 _17737_ (
    .A(_00061_),
    .B(_08007_),
    .X(_08008_)
  );
  sg13g2_o21ai_1 _17738_ (
    .A1(_08188_),
    .A2(_09502_),
    .B1(addr_i_5_),
    .Y(_08009_)
  );
  sg13g2_o21ai_1 _17739_ (
    .A1(_08188_),
    .A2(_00209_),
    .B1(addr_i_4_),
    .Y(_08010_)
  );
  sg13g2_a21oi_1 _17740_ (
    .A1(_08009_),
    .A2(_08010_),
    .B1(_04191_),
    .Y(_08012_)
  );
  sg13g2_a21oi_1 _17741_ (
    .A1(_03281_),
    .A2(_01966_),
    .B1(_01232_),
    .Y(_08013_)
  );
  sg13g2_o21ai_1 _17742_ (
    .A1(addr_i_4_),
    .A2(_08013_),
    .B1(_00907_),
    .Y(_08014_)
  );
  sg13g2_o21ai_1 _17743_ (
    .A1(_08012_),
    .A2(_08014_),
    .B1(addr_i_3_),
    .Y(_08015_)
  );
  sg13g2_o21ai_1 _17744_ (
    .A1(_00409_),
    .A2(_01499_),
    .B1(_08015_),
    .Y(_08016_)
  );
  sg13g2_o21ai_1 _17745_ (
    .A1(_08008_),
    .A2(_08016_),
    .B1(_00423_),
    .Y(_08017_)
  );
  sg13g2_o21ai_1 _17746_ (
    .A1(addr_i_5_),
    .A2(_07643_),
    .B1(_02002_),
    .Y(_08018_)
  );
  sg13g2_nand2_1 _17747_ (
    .A(_01946_),
    .B(_02546_),
    .Y(_08019_)
  );
  sg13g2_o21ai_1 _17748_ (
    .A1(addr_i_2_),
    .A2(_02152_),
    .B1(addr_i_3_),
    .Y(_08020_)
  );
  sg13g2_a21oi_1 _17749_ (
    .A1(_01353_),
    .A2(_08020_),
    .B1(_02064_),
    .Y(_08021_)
  );
  sg13g2_a22oi_1 _17750_ (
    .A1(addr_i_5_),
    .A2(_08019_),
    .B1(_08021_),
    .B2(_09183_),
    .Y(_08023_)
  );
  sg13g2_a21oi_1 _17751_ (
    .A1(_01339_),
    .A2(_04754_),
    .B1(_01543_),
    .Y(_08024_)
  );
  sg13g2_a22oi_1 _17752_ (
    .A1(_00993_),
    .A2(_01747_),
    .B1(_08024_),
    .B2(_00659_),
    .Y(_08025_)
  );
  sg13g2_a21oi_1 _17753_ (
    .A1(_08399_),
    .A2(_08023_),
    .B1(_08025_),
    .Y(_08026_)
  );
  sg13g2_a22oi_1 _17754_ (
    .A1(_09474_),
    .A2(_08018_),
    .B1(_08026_),
    .B2(_03259_),
    .Y(_08027_)
  );
  sg13g2_o21ai_1 _17755_ (
    .A1(addr_i_3_),
    .A2(_01057_),
    .B1(_05490_),
    .Y(_08028_)
  );
  sg13g2_a21oi_1 _17756_ (
    .A1(_05780_),
    .A2(_01050_),
    .B1(_00701_),
    .Y(_08029_)
  );
  sg13g2_a22oi_1 _17757_ (
    .A1(addr_i_5_),
    .A2(_08028_),
    .B1(_08029_),
    .B2(_01387_),
    .Y(_08030_)
  );
  sg13g2_and2_1 _17758_ (
    .A(_00391_),
    .B(_01305_),
    .X(_08031_)
  );
  sg13g2_a22oi_1 _17759_ (
    .A1(_00497_),
    .A2(_00712_),
    .B1(_03359_),
    .B2(_00899_),
    .Y(_08032_)
  );
  sg13g2_o21ai_1 _17760_ (
    .A1(_00051_),
    .A2(_00409_),
    .B1(_03617_),
    .Y(_08034_)
  );
  sg13g2_a22oi_1 _17761_ (
    .A1(_02641_),
    .A2(_08031_),
    .B1(_08032_),
    .B2(_08034_),
    .Y(_08035_)
  );
  sg13g2_o21ai_1 _17762_ (
    .A1(addr_i_7_),
    .A2(_08030_),
    .B1(_08035_),
    .Y(_08036_)
  );
  sg13g2_nand3b_1 _17763_ (
    .A_N(_08027_),
    .B(_08036_),
    .C(addr_i_9_),
    .Y(_08037_)
  );
  sg13g2_nand4_1 _17764_ (
    .A(addr_i_10_),
    .B(_08004_),
    .C(_08017_),
    .D(_08037_),
    .Y(_08038_)
  );
  sg13g2_o21ai_1 _17765_ (
    .A1(_01587_),
    .A2(_00597_),
    .B1(_02990_),
    .Y(_08039_)
  );
  sg13g2_o21ai_1 _17766_ (
    .A1(addr_i_7_),
    .A2(_03288_),
    .B1(_08653_),
    .Y(_08040_)
  );
  sg13g2_nand3_1 _17767_ (
    .A(_01499_),
    .B(_08039_),
    .C(_08040_),
    .Y(_08041_)
  );
  sg13g2_a21oi_1 _17768_ (
    .A1(_09510_),
    .A2(_01579_),
    .B1(_08188_),
    .Y(_08042_)
  );
  sg13g2_o21ai_1 _17769_ (
    .A1(addr_i_2_),
    .A2(_08042_),
    .B1(_09271_),
    .Y(_08043_)
  );
  sg13g2_o21ai_1 _17770_ (
    .A1(_00581_),
    .A2(_02623_),
    .B1(addr_i_3_),
    .Y(_08046_)
  );
  sg13g2_a22oi_1 _17771_ (
    .A1(_05811_),
    .A2(_06473_),
    .B1(_08046_),
    .B2(_01232_),
    .Y(_08047_)
  );
  sg13g2_nor3_1 _17772_ (
    .A(addr_i_3_),
    .B(_01292_),
    .C(_01627_),
    .Y(_08048_)
  );
  sg13g2_o21ai_1 _17773_ (
    .A1(_08047_),
    .A2(_08048_),
    .B1(addr_i_4_),
    .Y(_08049_)
  );
  sg13g2_o21ai_1 _17774_ (
    .A1(_08041_),
    .A2(_08043_),
    .B1(_08049_),
    .Y(_08050_)
  );
  sg13g2_a21o_1 _17775_ (
    .A1(_00884_),
    .A2(_03324_),
    .B1(addr_i_2_),
    .X(_08051_)
  );
  sg13g2_nand2_1 _17776_ (
    .A(_09513_),
    .B(_01398_),
    .Y(_08052_)
  );
  sg13g2_a22oi_1 _17777_ (
    .A1(addr_i_2_),
    .A2(_08052_),
    .B1(_00346_),
    .B2(_04672_),
    .Y(_08053_)
  );
  sg13g2_a21oi_1 _17778_ (
    .A1(_00441_),
    .A2(_06132_),
    .B1(_01970_),
    .Y(_08054_)
  );
  sg13g2_nor2_1 _17779_ (
    .A(_00200_),
    .B(_03962_),
    .Y(_08055_)
  );
  sg13g2_a21oi_1 _17780_ (
    .A1(_04162_),
    .A2(_01252_),
    .B1(addr_i_3_),
    .Y(_08057_)
  );
  sg13g2_nor4_1 _17781_ (
    .A(_07603_),
    .B(_08054_),
    .C(_08055_),
    .D(_08057_),
    .Y(_08058_)
  );
  sg13g2_o21ai_1 _17782_ (
    .A1(_00244_),
    .A2(_02424_),
    .B1(addr_i_3_),
    .Y(_08059_)
  );
  sg13g2_a21oi_1 _17783_ (
    .A1(_00651_),
    .A2(_08059_),
    .B1(_02179_),
    .Y(_08060_)
  );
  sg13g2_a22oi_1 _17784_ (
    .A1(_08051_),
    .A2(_08053_),
    .B1(_08058_),
    .B2(_08060_),
    .Y(_08061_)
  );
  sg13g2_o21ai_1 _17785_ (
    .A1(_01151_),
    .A2(_08050_),
    .B1(_08061_),
    .Y(_08062_)
  );
  sg13g2_nor3_1 _17786_ (
    .A(_00778_),
    .B(_00838_),
    .C(_04681_),
    .Y(_08063_)
  );
  sg13g2_a22oi_1 _17787_ (
    .A1(addr_i_3_),
    .A2(_05921_),
    .B1(_00667_),
    .B2(addr_i_7_),
    .Y(_08064_)
  );
  sg13g2_or3_1 _17788_ (
    .A(addr_i_5_),
    .B(_08063_),
    .C(_08064_),
    .X(_08065_)
  );
  sg13g2_a21oi_1 _17789_ (
    .A1(_00051_),
    .A2(_02467_),
    .B1(_02530_),
    .Y(_08066_)
  );
  sg13g2_a21oi_1 _17790_ (
    .A1(_00191_),
    .A2(_00449_),
    .B1(_08066_),
    .Y(_08068_)
  );
  sg13g2_o21ai_1 _17791_ (
    .A1(_02330_),
    .A2(_03433_),
    .B1(addr_i_4_),
    .Y(_08069_)
  );
  sg13g2_nand3_1 _17792_ (
    .A(_08065_),
    .B(_08068_),
    .C(_08069_),
    .Y(_08070_)
  );
  sg13g2_nand2_1 _17793_ (
    .A(addr_i_3_),
    .B(_02081_),
    .Y(_08071_)
  );
  sg13g2_o21ai_1 _17794_ (
    .A1(_01420_),
    .A2(_03267_),
    .B1(addr_i_5_),
    .Y(_08072_)
  );
  sg13g2_nand3_1 _17795_ (
    .A(_03361_),
    .B(_08071_),
    .C(_08072_),
    .Y(_08073_)
  );
  sg13g2_a21oi_1 _17796_ (
    .A1(_00573_),
    .A2(_00968_),
    .B1(addr_i_5_),
    .Y(_08074_)
  );
  sg13g2_a22oi_1 _17797_ (
    .A1(_00386_),
    .A2(_05220_),
    .B1(_08074_),
    .B2(addr_i_3_),
    .Y(_08075_)
  );
  sg13g2_nand2_1 _17798_ (
    .A(_00103_),
    .B(_02732_),
    .Y(_08076_)
  );
  sg13g2_a22oi_1 _17799_ (
    .A1(_00659_),
    .A2(_08076_),
    .B1(_05813_),
    .B2(_04754_),
    .Y(_08077_)
  );
  sg13g2_a22oi_1 _17800_ (
    .A1(_00818_),
    .A2(_02312_),
    .B1(_01611_),
    .B2(_01542_),
    .Y(_08079_)
  );
  sg13g2_o21ai_1 _17801_ (
    .A1(_08075_),
    .A2(_08077_),
    .B1(_08079_),
    .Y(_08080_)
  );
  sg13g2_nand3_1 _17802_ (
    .A(_01773_),
    .B(_08073_),
    .C(_08080_),
    .Y(_08081_)
  );
  sg13g2_a221oi_1 _17803_ (
    .A1(addr_i_9_),
    .A2(_08062_),
    .B1(_08070_),
    .B2(_00423_),
    .C1(_08081_),
    .Y(_08082_)
  );
  sg13g2_nor2_1 _17804_ (
    .A(_03051_),
    .B(_08082_),
    .Y(_08083_)
  );
  sg13g2_o21ai_1 _17805_ (
    .A1(addr_i_5_),
    .A2(_00375_),
    .B1(addr_i_2_),
    .Y(_08084_)
  );
  sg13g2_a21oi_1 _17806_ (
    .A1(_08084_),
    .A2(_03445_),
    .B1(_04672_),
    .Y(_08085_)
  );
  sg13g2_o21ai_1 _17807_ (
    .A1(_03012_),
    .A2(_02954_),
    .B1(_01224_),
    .Y(_08086_)
  );
  sg13g2_a21oi_1 _17808_ (
    .A1(_00148_),
    .A2(_03325_),
    .B1(_00951_),
    .Y(_08087_)
  );
  sg13g2_a21oi_1 _17809_ (
    .A1(addr_i_7_),
    .A2(_08086_),
    .B1(_08087_),
    .Y(_08088_)
  );
  sg13g2_a221oi_1 _17810_ (
    .A1(addr_i_7_),
    .A2(_03110_),
    .B1(_01745_),
    .B2(_00242_),
    .C1(_00354_),
    .Y(_08090_)
  );
  sg13g2_a22oi_1 _17811_ (
    .A1(_08388_),
    .A2(_02594_),
    .B1(_08090_),
    .B2(addr_i_2_),
    .Y(_08091_)
  );
  sg13g2_a21oi_1 _17812_ (
    .A1(_04572_),
    .A2(_01302_),
    .B1(_08091_),
    .Y(_08092_)
  );
  sg13g2_o21ai_1 _17813_ (
    .A1(_00146_),
    .A2(_08088_),
    .B1(_08092_),
    .Y(_08093_)
  );
  sg13g2_o21ai_1 _17814_ (
    .A1(_08863_),
    .A2(_03358_),
    .B1(_03660_),
    .Y(_08094_)
  );
  sg13g2_a21oi_1 _17815_ (
    .A1(addr_i_6_),
    .A2(_08094_),
    .B1(_06950_),
    .Y(_08095_)
  );
  sg13g2_o21ai_1 _17816_ (
    .A1(_00011_),
    .A2(_02153_),
    .B1(_08111_),
    .Y(_08096_)
  );
  sg13g2_o21ai_1 _17817_ (
    .A1(_07038_),
    .A2(_03324_),
    .B1(_08096_),
    .Y(_08097_)
  );
  sg13g2_nor2_1 _17818_ (
    .A(_00467_),
    .B(_01222_),
    .Y(_08098_)
  );
  sg13g2_a21oi_1 _17819_ (
    .A1(addr_i_2_),
    .A2(_08097_),
    .B1(_08098_),
    .Y(_08099_)
  );
  sg13g2_o21ai_1 _17820_ (
    .A1(addr_i_2_),
    .A2(_08095_),
    .B1(_08099_),
    .Y(_08101_)
  );
  sg13g2_mux2_1 _17821_ (
    .A0(_08093_),
    .A1(_08101_),
    .S(_00782_),
    .X(_08102_)
  );
  sg13g2_o21ai_1 _17822_ (
    .A1(_08085_),
    .A2(_08102_),
    .B1(addr_i_9_),
    .Y(_08103_)
  );
  sg13g2_nor3_1 _17823_ (
    .A(_00053_),
    .B(_00214_),
    .C(_00348_),
    .Y(_08104_)
  );
  sg13g2_o21ai_1 _17824_ (
    .A1(addr_i_4_),
    .A2(_01480_),
    .B1(addr_i_2_),
    .Y(_08105_)
  );
  sg13g2_a21oi_1 _17825_ (
    .A1(_04715_),
    .A2(_00284_),
    .B1(_01067_),
    .Y(_08106_)
  );
  sg13g2_o21ai_1 _17826_ (
    .A1(_02171_),
    .A2(_08106_),
    .B1(addr_i_4_),
    .Y(_08107_)
  );
  sg13g2_nor2_1 _17827_ (
    .A(_05457_),
    .B(_02462_),
    .Y(_08108_)
  );
  sg13g2_o21ai_1 _17828_ (
    .A1(_02750_),
    .A2(_08108_),
    .B1(_02063_),
    .Y(_08109_)
  );
  sg13g2_a21oi_1 _17829_ (
    .A1(_08107_),
    .A2(_08109_),
    .B1(_00588_),
    .Y(_08110_)
  );
  sg13g2_a21oi_1 _17830_ (
    .A1(_07724_),
    .A2(_09475_),
    .B1(addr_i_3_),
    .Y(_08112_)
  );
  sg13g2_o21ai_1 _17831_ (
    .A1(_09493_),
    .A2(_01014_),
    .B1(addr_i_3_),
    .Y(_08113_)
  );
  sg13g2_o21ai_1 _17832_ (
    .A1(addr_i_4_),
    .A2(_02583_),
    .B1(_08113_),
    .Y(_08114_)
  );
  sg13g2_o21ai_1 _17833_ (
    .A1(_08112_),
    .A2(_08114_),
    .B1(_07934_),
    .Y(_08115_)
  );
  sg13g2_nand3_1 _17834_ (
    .A(_01047_),
    .B(_01144_),
    .C(_02494_),
    .Y(_08116_)
  );
  sg13g2_nand3_1 _17835_ (
    .A(addr_i_10_),
    .B(_08115_),
    .C(_08116_),
    .Y(_08117_)
  );
  sg13g2_or2_1 _17836_ (
    .A(_08110_),
    .B(_08117_),
    .X(_08118_)
  );
  sg13g2_nand3_1 _17837_ (
    .A(_00573_),
    .B(_02607_),
    .C(_05334_),
    .Y(_08119_)
  );
  sg13g2_a221oi_1 _17838_ (
    .A1(_01336_),
    .A2(_05081_),
    .B1(_00862_),
    .B2(_00068_),
    .C1(_08119_),
    .Y(_08120_)
  );
  sg13g2_a221oi_1 _17839_ (
    .A1(_08104_),
    .A2(_08105_),
    .B1(_08118_),
    .B2(_02221_),
    .C1(_08120_),
    .Y(_08121_)
  );
  sg13g2_o21ai_1 _17840_ (
    .A1(_05999_),
    .A2(_02441_),
    .B1(addr_i_3_),
    .Y(_08123_)
  );
  sg13g2_o21ai_1 _17841_ (
    .A1(_00376_),
    .A2(_02792_),
    .B1(_03281_),
    .Y(_08124_)
  );
  sg13g2_nand3_1 _17842_ (
    .A(_01517_),
    .B(_08123_),
    .C(_08124_),
    .Y(_08125_)
  );
  sg13g2_o21ai_1 _17843_ (
    .A1(_02141_),
    .A2(_03864_),
    .B1(_03875_),
    .Y(_08126_)
  );
  sg13g2_a21oi_1 _17844_ (
    .A1(_00938_),
    .A2(_01432_),
    .B1(addr_i_4_),
    .Y(_08127_)
  );
  sg13g2_o21ai_1 _17845_ (
    .A1(addr_i_3_),
    .A2(_00687_),
    .B1(addr_i_7_),
    .Y(_08128_)
  );
  sg13g2_a22oi_1 _17846_ (
    .A1(addr_i_4_),
    .A2(_08126_),
    .B1(_08127_),
    .B2(_08128_),
    .Y(_08129_)
  );
  sg13g2_nor2_1 _17847_ (
    .A(_07282_),
    .B(_08129_),
    .Y(_08130_)
  );
  sg13g2_a221oi_1 _17848_ (
    .A1(_03270_),
    .A2(_07237_),
    .B1(_00304_),
    .B2(_00117_),
    .C1(_05856_),
    .Y(_08131_)
  );
  sg13g2_nand3_1 _17849_ (
    .A(_00347_),
    .B(_01589_),
    .C(_09415_),
    .Y(_08132_)
  );
  sg13g2_nand2b_1 _17850_ (
    .A_N(_08131_),
    .B(_08132_),
    .Y(_08134_)
  );
  sg13g2_nor3_1 _17851_ (
    .A(addr_i_3_),
    .B(_07967_),
    .C(_00304_),
    .Y(_08135_)
  );
  sg13g2_o21ai_1 _17852_ (
    .A1(_01590_),
    .A2(_08135_),
    .B1(addr_i_5_),
    .Y(_08136_)
  );
  sg13g2_a21oi_1 _17853_ (
    .A1(_08134_),
    .A2(_08136_),
    .B1(_01099_),
    .Y(_08137_)
  );
  sg13g2_a21oi_1 _17854_ (
    .A1(_01432_),
    .A2(_06324_),
    .B1(addr_i_4_),
    .Y(_08138_)
  );
  sg13g2_a21oi_1 _17855_ (
    .A1(_09510_),
    .A2(_00831_),
    .B1(_01674_),
    .Y(_08139_)
  );
  sg13g2_a21oi_1 _17856_ (
    .A1(_00482_),
    .A2(_05780_),
    .B1(addr_i_3_),
    .Y(_08140_)
  );
  sg13g2_nor4_1 _17857_ (
    .A(_07603_),
    .B(_08138_),
    .C(_08139_),
    .D(_08140_),
    .Y(_08141_)
  );
  sg13g2_a22oi_1 _17858_ (
    .A1(_08125_),
    .A2(_08130_),
    .B1(_08137_),
    .B2(_08141_),
    .Y(_08142_)
  );
  sg13g2_or2_1 _17859_ (
    .A(_03776_),
    .B(_03061_),
    .X(_08143_)
  );
  sg13g2_o21ai_1 _17860_ (
    .A1(_06795_),
    .A2(_05568_),
    .B1(_00999_),
    .Y(_08145_)
  );
  sg13g2_o21ai_1 _17861_ (
    .A1(_00060_),
    .A2(_08143_),
    .B1(_08145_),
    .Y(_08146_)
  );
  sg13g2_or2_1 _17862_ (
    .A(_04041_),
    .B(_01305_),
    .X(_08147_)
  );
  sg13g2_nor3_1 _17863_ (
    .A(_00115_),
    .B(_06010_),
    .C(_02443_),
    .Y(_08148_)
  );
  sg13g2_a22oi_1 _17864_ (
    .A1(_00701_),
    .A2(_08147_),
    .B1(_08148_),
    .B2(_01099_),
    .Y(_08149_)
  );
  sg13g2_a22oi_1 _17865_ (
    .A1(_00708_),
    .A2(_08146_),
    .B1(_08149_),
    .B2(addr_i_9_),
    .Y(_08150_)
  );
  sg13g2_a21oi_1 _17866_ (
    .A1(addr_i_9_),
    .A2(_08142_),
    .B1(_08150_),
    .Y(_08151_)
  );
  sg13g2_nand2_1 _17867_ (
    .A(addr_i_5_),
    .B(_02076_),
    .Y(_08152_)
  );
  sg13g2_a22oi_1 _17868_ (
    .A1(_06717_),
    .A2(_08152_),
    .B1(_00285_),
    .B2(_02277_),
    .Y(_08153_)
  );
  sg13g2_nor2_1 _17869_ (
    .A(_04225_),
    .B(_08153_),
    .Y(_08154_)
  );
  sg13g2_nor2_1 _17870_ (
    .A(_05723_),
    .B(_08154_),
    .Y(_08157_)
  );
  sg13g2_nor2_1 _17871_ (
    .A(_02963_),
    .B(_08157_),
    .Y(_08158_)
  );
  sg13g2_nor3_1 _17872_ (
    .A(_03497_),
    .B(_09260_),
    .C(_03494_),
    .Y(_08159_)
  );
  sg13g2_nor4_1 _17873_ (
    .A(addr_i_10_),
    .B(_08151_),
    .C(_08158_),
    .D(_08159_),
    .Y(_08160_)
  );
  sg13g2_a22oi_1 _17874_ (
    .A1(_08103_),
    .A2(_08121_),
    .B1(_08160_),
    .B2(addr_i_11_),
    .Y(_08161_)
  );
  sg13g2_a22oi_1 _17875_ (
    .A1(_08038_),
    .A2(_08083_),
    .B1(_08161_),
    .B2(addr_i_12_),
    .Y(_08162_)
  );
  sg13g2_a21oi_1 _17876_ (
    .A1(addr_i_12_),
    .A2(_07991_),
    .B1(_08162_),
    .Y(data_o_4_)
  );
  sg13g2_o21ai_1 _17877_ (
    .A1(_02542_),
    .A2(_03562_),
    .B1(_00048_),
    .Y(_08163_)
  );
  sg13g2_a21oi_1 _17878_ (
    .A1(_04442_),
    .A2(_02772_),
    .B1(_05834_),
    .Y(_08164_)
  );
  sg13g2_nand2_1 _17879_ (
    .A(_08163_),
    .B(_08164_),
    .Y(_08165_)
  );
  sg13g2_a21oi_1 _17880_ (
    .A1(_00500_),
    .A2(_07427_),
    .B1(_03631_),
    .Y(_08167_)
  );
  sg13g2_a21oi_1 _17881_ (
    .A1(_09492_),
    .A2(_03288_),
    .B1(_02428_),
    .Y(_08168_)
  );
  sg13g2_o21ai_1 _17882_ (
    .A1(_00747_),
    .A2(_08168_),
    .B1(_06695_),
    .Y(_08169_)
  );
  sg13g2_nand2_1 _17883_ (
    .A(_06088_),
    .B(_02405_),
    .Y(_08170_)
  );
  sg13g2_a22oi_1 _17884_ (
    .A1(_00967_),
    .A2(_08170_),
    .B1(_02632_),
    .B2(_00060_),
    .Y(_08171_)
  );
  sg13g2_o21ai_1 _17885_ (
    .A1(addr_i_3_),
    .A2(_00842_),
    .B1(_04191_),
    .Y(_08172_)
  );
  sg13g2_nor2_1 _17886_ (
    .A(_08171_),
    .B(_08172_),
    .Y(_08173_)
  );
  sg13g2_nor2_1 _17887_ (
    .A(_08169_),
    .B(_08173_),
    .Y(_08174_)
  );
  sg13g2_a22oi_1 _17888_ (
    .A1(addr_i_8_),
    .A2(_08167_),
    .B1(_08174_),
    .B2(addr_i_9_),
    .Y(_08175_)
  );
  sg13g2_a21oi_1 _17889_ (
    .A1(addr_i_9_),
    .A2(_04606_),
    .B1(_08175_),
    .Y(_08176_)
  );
  sg13g2_nor2_1 _17890_ (
    .A(addr_i_10_),
    .B(_08176_),
    .Y(_08178_)
  );
  sg13g2_a22oi_1 _17891_ (
    .A1(_01646_),
    .A2(_08165_),
    .B1(_08178_),
    .B2(_01359_),
    .Y(_08179_)
  );
  sg13g2_nor2_1 _17892_ (
    .A(_06143_),
    .B(_01276_),
    .Y(_08180_)
  );
  sg13g2_a21oi_1 _17893_ (
    .A1(addr_i_4_),
    .A2(_08180_),
    .B1(_02424_),
    .Y(_08181_)
  );
  sg13g2_nor2_1 _17894_ (
    .A(_06619_),
    .B(_08181_),
    .Y(_08182_)
  );
  sg13g2_a21oi_1 _17895_ (
    .A1(_00500_),
    .A2(_02091_),
    .B1(_08182_),
    .Y(_08183_)
  );
  sg13g2_nand2_1 _17896_ (
    .A(_02694_),
    .B(_01791_),
    .Y(_08184_)
  );
  sg13g2_a21oi_1 _17897_ (
    .A1(_01729_),
    .A2(_04371_),
    .B1(addr_i_7_),
    .Y(_08185_)
  );
  sg13g2_a22oi_1 _17898_ (
    .A1(addr_i_4_),
    .A2(_08184_),
    .B1(_08185_),
    .B2(addr_i_3_),
    .Y(_08186_)
  );
  sg13g2_a21oi_1 _17899_ (
    .A1(addr_i_3_),
    .A2(_08183_),
    .B1(_08186_),
    .Y(_08187_)
  );
  sg13g2_nand2_1 _17900_ (
    .A(addr_i_8_),
    .B(_02738_),
    .Y(_08189_)
  );
  sg13g2_o21ai_1 _17901_ (
    .A1(addr_i_4_),
    .A2(_01212_),
    .B1(_02165_),
    .Y(_08190_)
  );
  sg13g2_a21oi_1 _17902_ (
    .A1(addr_i_2_),
    .A2(_03964_),
    .B1(_00467_),
    .Y(_08191_)
  );
  sg13g2_a22oi_1 _17903_ (
    .A1(addr_i_3_),
    .A2(_08190_),
    .B1(_08191_),
    .B2(_04778_),
    .Y(_08192_)
  );
  sg13g2_nor2_1 _17904_ (
    .A(_08056_),
    .B(_00951_),
    .Y(_08193_)
  );
  sg13g2_a21oi_1 _17905_ (
    .A1(_00315_),
    .A2(_01230_),
    .B1(_00070_),
    .Y(_08194_)
  );
  sg13g2_a22oi_1 _17906_ (
    .A1(_02858_),
    .A2(_08193_),
    .B1(_08194_),
    .B2(addr_i_8_),
    .Y(_08195_)
  );
  sg13g2_o21ai_1 _17907_ (
    .A1(addr_i_6_),
    .A2(_08192_),
    .B1(_08195_),
    .Y(_08196_)
  );
  sg13g2_o21ai_1 _17908_ (
    .A1(_08187_),
    .A2(_08189_),
    .B1(_08196_),
    .Y(_08197_)
  );
  sg13g2_a21oi_1 _17909_ (
    .A1(_00505_),
    .A2(_05501_),
    .B1(_02632_),
    .Y(_08198_)
  );
  sg13g2_a22oi_1 _17910_ (
    .A1(_09061_),
    .A2(_00226_),
    .B1(_01977_),
    .B2(_03589_),
    .Y(_08200_)
  );
  sg13g2_o21ai_1 _17911_ (
    .A1(addr_i_5_),
    .A2(_08198_),
    .B1(_08200_),
    .Y(_08201_)
  );
  sg13g2_o21ai_1 _17912_ (
    .A1(_02191_),
    .A2(_04328_),
    .B1(addr_i_8_),
    .Y(_08202_)
  );
  sg13g2_nor3_1 _17913_ (
    .A(_02343_),
    .B(addr_i_5_),
    .C(_02426_),
    .Y(_08203_)
  );
  sg13g2_o21ai_1 _17914_ (
    .A1(_00087_),
    .A2(_08203_),
    .B1(addr_i_4_),
    .Y(_08204_)
  );
  sg13g2_nor2_1 _17915_ (
    .A(addr_i_4_),
    .B(_07769_),
    .Y(_08205_)
  );
  sg13g2_a21oi_1 _17916_ (
    .A1(addr_i_6_),
    .A2(_00090_),
    .B1(_08205_),
    .Y(_08206_)
  );
  sg13g2_a21oi_1 _17917_ (
    .A1(_08204_),
    .A2(_08206_),
    .B1(addr_i_3_),
    .Y(_08207_)
  );
  sg13g2_a22oi_1 _17918_ (
    .A1(addr_i_3_),
    .A2(_08201_),
    .B1(_08202_),
    .B2(_08207_),
    .Y(_08208_)
  );
  sg13g2_a21oi_1 _17919_ (
    .A1(addr_i_3_),
    .A2(_08376_),
    .B1(_00738_),
    .Y(_08209_)
  );
  sg13g2_o21ai_1 _17920_ (
    .A1(addr_i_6_),
    .A2(_08209_),
    .B1(_01060_),
    .Y(_08211_)
  );
  sg13g2_a21oi_1 _17921_ (
    .A1(_00404_),
    .A2(_00985_),
    .B1(addr_i_4_),
    .Y(_08212_)
  );
  sg13g2_o21ai_1 _17922_ (
    .A1(_01308_),
    .A2(_08211_),
    .B1(_08212_),
    .Y(_08213_)
  );
  sg13g2_a21oi_1 _17923_ (
    .A1(_01353_),
    .A2(_00603_),
    .B1(_08332_),
    .Y(_08214_)
  );
  sg13g2_o21ai_1 _17924_ (
    .A1(_00301_),
    .A2(_08214_),
    .B1(addr_i_4_),
    .Y(_08215_)
  );
  sg13g2_and4_1 _17925_ (
    .A(_03617_),
    .B(_03707_),
    .C(_08213_),
    .D(_08215_),
    .X(_08216_)
  );
  sg13g2_or3_1 _17926_ (
    .A(_01351_),
    .B(_08208_),
    .C(_08216_),
    .X(_08217_)
  );
  sg13g2_o21ai_1 _17927_ (
    .A1(addr_i_9_),
    .A2(_08197_),
    .B1(_08217_),
    .Y(_08218_)
  );
  sg13g2_o21ai_1 _17928_ (
    .A1(_02772_),
    .A2(_03980_),
    .B1(addr_i_3_),
    .Y(_08219_)
  );
  sg13g2_a22oi_1 _17929_ (
    .A1(_00061_),
    .A2(_00426_),
    .B1(_02273_),
    .B2(_01365_),
    .Y(_08220_)
  );
  sg13g2_o21ai_1 _17930_ (
    .A1(_00268_),
    .A2(_00159_),
    .B1(addr_i_3_),
    .Y(_08222_)
  );
  sg13g2_nand3_1 _17931_ (
    .A(_00440_),
    .B(_01983_),
    .C(_08222_),
    .Y(_08223_)
  );
  sg13g2_nor2_1 _17932_ (
    .A(_00517_),
    .B(_08223_),
    .Y(_08224_)
  );
  sg13g2_o21ai_1 _17933_ (
    .A1(addr_i_3_),
    .A2(_00275_),
    .B1(_00007_),
    .Y(_08225_)
  );
  sg13g2_a21oi_1 _17934_ (
    .A1(_04191_),
    .A2(_08225_),
    .B1(_00898_),
    .Y(_08226_)
  );
  sg13g2_nor2_1 _17935_ (
    .A(addr_i_4_),
    .B(_08226_),
    .Y(_08227_)
  );
  sg13g2_o21ai_1 _17936_ (
    .A1(addr_i_4_),
    .A2(_01972_),
    .B1(_09149_),
    .Y(_08228_)
  );
  sg13g2_a221oi_1 _17937_ (
    .A1(_06419_),
    .A2(_01603_),
    .B1(_07270_),
    .B2(_01441_),
    .C1(_08155_),
    .Y(_08229_)
  );
  sg13g2_a21oi_1 _17938_ (
    .A1(addr_i_2_),
    .A2(_08228_),
    .B1(_08229_),
    .Y(_08230_)
  );
  sg13g2_a21o_1 _17939_ (
    .A1(_01265_),
    .A2(_05464_),
    .B1(addr_i_7_),
    .X(_08231_)
  );
  sg13g2_o21ai_1 _17940_ (
    .A1(addr_i_6_),
    .A2(_08230_),
    .B1(_08231_),
    .Y(_08233_)
  );
  sg13g2_nor4_1 _17941_ (
    .A(_01151_),
    .B(_02772_),
    .C(_08227_),
    .D(_08233_),
    .Y(_08234_)
  );
  sg13g2_a22oi_1 _17942_ (
    .A1(_08219_),
    .A2(_08220_),
    .B1(_08224_),
    .B2(_08234_),
    .Y(_08235_)
  );
  sg13g2_a21oi_1 _17943_ (
    .A1(_04413_),
    .A2(_02956_),
    .B1(addr_i_7_),
    .Y(_08236_)
  );
  sg13g2_a21o_1 _17944_ (
    .A1(_00884_),
    .A2(_02002_),
    .B1(addr_i_6_),
    .X(_08237_)
  );
  sg13g2_o21ai_1 _17945_ (
    .A1(_00334_),
    .A2(_07064_),
    .B1(addr_i_4_),
    .Y(_08238_)
  );
  sg13g2_a21oi_1 _17946_ (
    .A1(_08237_),
    .A2(_08238_),
    .B1(_05822_),
    .Y(_08239_)
  );
  sg13g2_a22oi_1 _17947_ (
    .A1(_00073_),
    .A2(_01837_),
    .B1(_08236_),
    .B2(_08239_),
    .Y(_08240_)
  );
  sg13g2_nor2_1 _17948_ (
    .A(_08056_),
    .B(_02026_),
    .Y(_08241_)
  );
  sg13g2_o21ai_1 _17949_ (
    .A1(_00091_),
    .A2(_07248_),
    .B1(_00594_),
    .Y(_08242_)
  );
  sg13g2_o21ai_1 _17950_ (
    .A1(addr_i_6_),
    .A2(_08241_),
    .B1(_08242_),
    .Y(_08244_)
  );
  sg13g2_a21oi_1 _17951_ (
    .A1(_00034_),
    .A2(_03391_),
    .B1(addr_i_2_),
    .Y(_08245_)
  );
  sg13g2_o21ai_1 _17952_ (
    .A1(_08951_),
    .A2(_04655_),
    .B1(_04662_),
    .Y(_08246_)
  );
  sg13g2_nor4_1 _17953_ (
    .A(_03227_),
    .B(_00732_),
    .C(_08245_),
    .D(_08246_),
    .Y(_08247_)
  );
  sg13g2_a21oi_1 _17954_ (
    .A1(_00708_),
    .A2(_08244_),
    .B1(_08247_),
    .Y(_08248_)
  );
  sg13g2_o21ai_1 _17955_ (
    .A1(addr_i_8_),
    .A2(_08240_),
    .B1(_08248_),
    .Y(_08249_)
  );
  sg13g2_a21oi_1 _17956_ (
    .A1(_05214_),
    .A2(_08249_),
    .B1(_00513_),
    .Y(_08250_)
  );
  sg13g2_o21ai_1 _17957_ (
    .A1(_01211_),
    .A2(_08235_),
    .B1(_08250_),
    .Y(_08251_)
  );
  sg13g2_a21oi_1 _17958_ (
    .A1(_01774_),
    .A2(_08218_),
    .B1(_08251_),
    .Y(_08252_)
  );
  sg13g2_o21ai_1 _17959_ (
    .A1(_00401_),
    .A2(_00346_),
    .B1(addr_i_2_),
    .Y(_08253_)
  );
  sg13g2_nand2_1 _17960_ (
    .A(_01182_),
    .B(_08253_),
    .Y(_08255_)
  );
  sg13g2_nor2_1 _17961_ (
    .A(_00507_),
    .B(_06860_),
    .Y(_08256_)
  );
  sg13g2_a22oi_1 _17962_ (
    .A1(_00169_),
    .A2(_08255_),
    .B1(_08256_),
    .B2(_01612_),
    .Y(_08257_)
  );
  sg13g2_nor2_1 _17963_ (
    .A(_04097_),
    .B(_02513_),
    .Y(_08258_)
  );
  sg13g2_o21ai_1 _17964_ (
    .A1(_07889_),
    .A2(_02490_),
    .B1(addr_i_2_),
    .Y(_08259_)
  );
  sg13g2_a21oi_1 _17965_ (
    .A1(_01182_),
    .A2(_08259_),
    .B1(_00172_),
    .Y(_08260_)
  );
  sg13g2_o21ai_1 _17966_ (
    .A1(_08258_),
    .A2(_08260_),
    .B1(_05834_),
    .Y(_08261_)
  );
  sg13g2_o21ai_1 _17967_ (
    .A1(addr_i_6_),
    .A2(_01571_),
    .B1(_03964_),
    .Y(_08262_)
  );
  sg13g2_a21oi_1 _17968_ (
    .A1(_03424_),
    .A2(_00138_),
    .B1(addr_i_3_),
    .Y(_08263_)
  );
  sg13g2_a22oi_1 _17969_ (
    .A1(addr_i_2_),
    .A2(_08262_),
    .B1(_08263_),
    .B2(addr_i_4_),
    .Y(_08264_)
  );
  sg13g2_nor2_1 _17970_ (
    .A(addr_i_7_),
    .B(_04097_),
    .Y(_08267_)
  );
  sg13g2_a22oi_1 _17971_ (
    .A1(_00626_),
    .A2(_01673_),
    .B1(_08267_),
    .B2(_00084_),
    .Y(_08268_)
  );
  sg13g2_nor2_1 _17972_ (
    .A(_08264_),
    .B(_08268_),
    .Y(_08269_)
  );
  sg13g2_a21oi_1 _17973_ (
    .A1(_00434_),
    .A2(_01499_),
    .B1(_00048_),
    .Y(_08270_)
  );
  sg13g2_nor4_1 _17974_ (
    .A(_00029_),
    .B(_02368_),
    .C(_08269_),
    .D(_08270_),
    .Y(_08271_)
  );
  sg13g2_a22oi_1 _17975_ (
    .A1(_08257_),
    .A2(_08261_),
    .B1(_08271_),
    .B2(addr_i_10_),
    .Y(_08272_)
  );
  sg13g2_o21ai_1 _17976_ (
    .A1(_01542_),
    .A2(_00132_),
    .B1(addr_i_3_),
    .Y(_08273_)
  );
  sg13g2_o21ai_1 _17977_ (
    .A1(_01103_),
    .A2(_00194_),
    .B1(_08273_),
    .Y(_08274_)
  );
  sg13g2_o21ai_1 _17978_ (
    .A1(_03690_),
    .A2(_00940_),
    .B1(_03064_),
    .Y(_08275_)
  );
  sg13g2_nand2_1 _17979_ (
    .A(_00427_),
    .B(_01684_),
    .Y(_08276_)
  );
  sg13g2_a21oi_1 _17980_ (
    .A1(_04396_),
    .A2(_02675_),
    .B1(_02803_),
    .Y(_08278_)
  );
  sg13g2_a22oi_1 _17981_ (
    .A1(addr_i_3_),
    .A2(_08276_),
    .B1(_08278_),
    .B2(_00436_),
    .Y(_08279_)
  );
  sg13g2_nor2_1 _17982_ (
    .A(addr_i_5_),
    .B(_08279_),
    .Y(_08280_)
  );
  sg13g2_a22oi_1 _17983_ (
    .A1(_00015_),
    .A2(_08274_),
    .B1(_08275_),
    .B2(_08280_),
    .Y(_08281_)
  );
  sg13g2_a21oi_1 _17984_ (
    .A1(_07625_),
    .A2(_03108_),
    .B1(_00951_),
    .Y(_08282_)
  );
  sg13g2_o21ai_1 _17985_ (
    .A1(_03455_),
    .A2(_00305_),
    .B1(addr_i_3_),
    .Y(_08283_)
  );
  sg13g2_a21oi_1 _17986_ (
    .A1(_02187_),
    .A2(_08283_),
    .B1(_06630_),
    .Y(_08284_)
  );
  sg13g2_a221oi_1 _17987_ (
    .A1(_09138_),
    .A2(_02742_),
    .B1(_05231_),
    .B2(_07149_),
    .C1(addr_i_4_),
    .Y(_08285_)
  );
  sg13g2_a22oi_1 _17988_ (
    .A1(addr_i_4_),
    .A2(_04328_),
    .B1(_08285_),
    .B2(_00068_),
    .Y(_08286_)
  );
  sg13g2_nor4_1 _17989_ (
    .A(_06706_),
    .B(_08282_),
    .C(_08284_),
    .D(_08286_),
    .Y(_08287_)
  );
  sg13g2_o21ai_1 _17990_ (
    .A1(_08281_),
    .A2(_08287_),
    .B1(addr_i_9_),
    .Y(_08289_)
  );
  sg13g2_o21ai_1 _17991_ (
    .A1(_00069_),
    .A2(_03497_),
    .B1(_02546_),
    .Y(_08290_)
  );
  sg13g2_nand2_1 _17992_ (
    .A(_08785_),
    .B(_00275_),
    .Y(_08291_)
  );
  sg13g2_o21ai_1 _17993_ (
    .A1(_02271_),
    .A2(_01718_),
    .B1(_08291_),
    .Y(_08292_)
  );
  sg13g2_a21oi_1 _17994_ (
    .A1(addr_i_4_),
    .A2(_08292_),
    .B1(_02215_),
    .Y(_08293_)
  );
  sg13g2_nor2_1 _17995_ (
    .A(addr_i_2_),
    .B(_08293_),
    .Y(_08294_)
  );
  sg13g2_o21ai_1 _17996_ (
    .A1(_00317_),
    .A2(_01007_),
    .B1(_02759_),
    .Y(_08295_)
  );
  sg13g2_a21oi_1 _17997_ (
    .A1(_01729_),
    .A2(_00185_),
    .B1(addr_i_3_),
    .Y(_08296_)
  );
  sg13g2_a22oi_1 _17998_ (
    .A1(addr_i_2_),
    .A2(_08295_),
    .B1(_08296_),
    .B2(_00898_),
    .Y(_08297_)
  );
  sg13g2_nor2_1 _17999_ (
    .A(addr_i_4_),
    .B(_08297_),
    .Y(_08298_)
  );
  sg13g2_a22oi_1 _18000_ (
    .A1(addr_i_2_),
    .A2(_08290_),
    .B1(_08294_),
    .B2(_08298_),
    .Y(_08300_)
  );
  sg13g2_a21oi_1 _18001_ (
    .A1(_02528_),
    .A2(_01343_),
    .B1(addr_i_4_),
    .Y(_08301_)
  );
  sg13g2_a221oi_1 _18002_ (
    .A1(addr_i_4_),
    .A2(_02437_),
    .B1(_02980_),
    .B2(addr_i_2_),
    .C1(_08301_),
    .Y(_08302_)
  );
  sg13g2_inv_1 _18003_ (
    .A(_08302_),
    .Y(_08303_)
  );
  sg13g2_nor2_1 _18004_ (
    .A(addr_i_4_),
    .B(_01587_),
    .Y(_08304_)
  );
  sg13g2_a22oi_1 _18005_ (
    .A1(addr_i_2_),
    .A2(_07744_),
    .B1(_07583_),
    .B2(_08304_),
    .Y(_08305_)
  );
  sg13g2_nand2b_1 _18006_ (
    .A_N(_08305_),
    .B(addr_i_6_),
    .Y(_08306_)
  );
  sg13g2_o21ai_1 _18007_ (
    .A1(_01587_),
    .A2(_02513_),
    .B1(_01070_),
    .Y(_08307_)
  );
  sg13g2_a21oi_1 _18008_ (
    .A1(_03930_),
    .A2(_08307_),
    .B1(_09359_),
    .Y(_08308_)
  );
  sg13g2_a21oi_1 _18009_ (
    .A1(_08306_),
    .A2(_08308_),
    .B1(addr_i_3_),
    .Y(_08309_)
  );
  sg13g2_a22oi_1 _18010_ (
    .A1(addr_i_3_),
    .A2(_08303_),
    .B1(_08309_),
    .B2(_04281_),
    .Y(_08311_)
  );
  sg13g2_nor2_1 _18011_ (
    .A(addr_i_8_),
    .B(_08311_),
    .Y(_08312_)
  );
  sg13g2_a22oi_1 _18012_ (
    .A1(addr_i_8_),
    .A2(_08300_),
    .B1(_08312_),
    .B2(_00109_),
    .Y(_08313_)
  );
  sg13g2_nand2_1 _18013_ (
    .A(_09483_),
    .B(_03195_),
    .Y(_08314_)
  );
  sg13g2_a22oi_1 _18014_ (
    .A1(_00191_),
    .A2(_08314_),
    .B1(_00850_),
    .B2(_09359_),
    .Y(_08315_)
  );
  sg13g2_a21oi_1 _18015_ (
    .A1(_00747_),
    .A2(_02746_),
    .B1(_01481_),
    .Y(_08316_)
  );
  sg13g2_a22oi_1 _18016_ (
    .A1(_04022_),
    .A2(_02652_),
    .B1(_08316_),
    .B2(addr_i_8_),
    .Y(_08317_)
  );
  sg13g2_o21ai_1 _18017_ (
    .A1(_05834_),
    .A2(_08315_),
    .B1(_08317_),
    .Y(_08318_)
  );
  sg13g2_nand4_1 _18018_ (
    .A(_09487_),
    .B(_00409_),
    .C(_05517_),
    .D(_05569_),
    .Y(_08319_)
  );
  sg13g2_nand2_1 _18019_ (
    .A(_00022_),
    .B(_01216_),
    .Y(_08320_)
  );
  sg13g2_nor2_1 _18020_ (
    .A(addr_i_3_),
    .B(_04355_),
    .Y(_08322_)
  );
  sg13g2_nor2_1 _18021_ (
    .A(_01114_),
    .B(_08609_),
    .Y(_08323_)
  );
  sg13g2_nor2_1 _18022_ (
    .A(_08322_),
    .B(_08323_),
    .Y(_08324_)
  );
  sg13g2_nand4_1 _18023_ (
    .A(addr_i_7_),
    .B(_08320_),
    .C(_08222_),
    .D(_08324_),
    .Y(_08325_)
  );
  sg13g2_nand3_1 _18024_ (
    .A(addr_i_4_),
    .B(_07337_),
    .C(_00315_),
    .Y(_08326_)
  );
  sg13g2_nand3_1 _18025_ (
    .A(_09474_),
    .B(_06909_),
    .C(_08326_),
    .Y(_08327_)
  );
  sg13g2_nand4_1 _18026_ (
    .A(addr_i_8_),
    .B(_08319_),
    .C(_08325_),
    .D(_08327_),
    .Y(_08328_)
  );
  sg13g2_nand3_1 _18027_ (
    .A(_01176_),
    .B(_08318_),
    .C(_08328_),
    .Y(_08329_)
  );
  sg13g2_nand2b_1 _18028_ (
    .A_N(_01451_),
    .B(_08329_),
    .Y(_08330_)
  );
  sg13g2_a22oi_1 _18029_ (
    .A1(_08272_),
    .A2(_08289_),
    .B1(_08313_),
    .B2(_08330_),
    .Y(_08331_)
  );
  sg13g2_o21ai_1 _18030_ (
    .A1(_03765_),
    .A2(_01917_),
    .B1(addr_i_2_),
    .Y(_08333_)
  );
  sg13g2_a21oi_1 _18031_ (
    .A1(_05116_),
    .A2(_08333_),
    .B1(addr_i_3_),
    .Y(_08334_)
  );
  sg13g2_nand2_1 _18032_ (
    .A(addr_i_3_),
    .B(_00447_),
    .Y(_08335_)
  );
  sg13g2_a21oi_1 _18033_ (
    .A1(_06310_),
    .A2(_08335_),
    .B1(_08696_),
    .Y(_08336_)
  );
  sg13g2_nor2_1 _18034_ (
    .A(_08334_),
    .B(_08336_),
    .Y(_08337_)
  );
  sg13g2_o21ai_1 _18035_ (
    .A1(_02470_),
    .A2(_01933_),
    .B1(_08337_),
    .Y(_08338_)
  );
  sg13g2_nor3_1 _18036_ (
    .A(_02732_),
    .B(_06198_),
    .C(_05112_),
    .Y(_08339_)
  );
  sg13g2_o21ai_1 _18037_ (
    .A1(addr_i_8_),
    .A2(_06099_),
    .B1(_02107_),
    .Y(_08340_)
  );
  sg13g2_a21oi_1 _18038_ (
    .A1(_06331_),
    .A2(_00943_),
    .B1(_05102_),
    .Y(_08341_)
  );
  sg13g2_a21oi_1 _18039_ (
    .A1(_08340_),
    .A2(_08341_),
    .B1(addr_i_4_),
    .Y(_08342_)
  );
  sg13g2_a22oi_1 _18040_ (
    .A1(addr_i_4_),
    .A2(_08338_),
    .B1(_08339_),
    .B2(_08342_),
    .Y(_08344_)
  );
  sg13g2_o21ai_1 _18041_ (
    .A1(addr_i_4_),
    .A2(_05902_),
    .B1(_05898_),
    .Y(_08345_)
  );
  sg13g2_a21oi_1 _18042_ (
    .A1(_00571_),
    .A2(_00940_),
    .B1(addr_i_8_),
    .Y(_08346_)
  );
  sg13g2_a21o_1 _18043_ (
    .A1(addr_i_3_),
    .A2(_08345_),
    .B1(_08346_),
    .X(_08347_)
  );
  sg13g2_nand3_1 _18044_ (
    .A(addr_i_8_),
    .B(_00238_),
    .C(_05910_),
    .Y(_08348_)
  );
  sg13g2_or3_1 _18045_ (
    .A(addr_i_2_),
    .B(addr_i_8_),
    .C(addr_i_6_),
    .X(_08349_)
  );
  sg13g2_a21oi_1 _18046_ (
    .A1(_01965_),
    .A2(_08349_),
    .B1(addr_i_3_),
    .Y(_08350_)
  );
  sg13g2_nor2_1 _18047_ (
    .A(_02459_),
    .B(_02780_),
    .Y(_08351_)
  );
  sg13g2_o21ai_1 _18048_ (
    .A1(_08350_),
    .A2(_08351_),
    .B1(_00354_),
    .Y(_08352_)
  );
  sg13g2_a21oi_1 _18049_ (
    .A1(_08348_),
    .A2(_08352_),
    .B1(addr_i_5_),
    .Y(_08353_)
  );
  sg13g2_a221oi_1 _18050_ (
    .A1(_01500_),
    .A2(_00156_),
    .B1(_08347_),
    .B2(addr_i_5_),
    .C1(_08353_),
    .Y(_08355_)
  );
  sg13g2_nor2_1 _18051_ (
    .A(addr_i_7_),
    .B(_08355_),
    .Y(_08356_)
  );
  sg13g2_a21oi_1 _18052_ (
    .A1(addr_i_7_),
    .A2(_08344_),
    .B1(_08356_),
    .Y(_08357_)
  );
  sg13g2_a21oi_1 _18053_ (
    .A1(_02696_),
    .A2(_05012_),
    .B1(addr_i_7_),
    .Y(_08358_)
  );
  sg13g2_a22oi_1 _18054_ (
    .A1(addr_i_7_),
    .A2(_03299_),
    .B1(_08358_),
    .B2(_00192_),
    .Y(_08359_)
  );
  sg13g2_nand3_1 _18055_ (
    .A(_00016_),
    .B(_01273_),
    .C(_01954_),
    .Y(_08360_)
  );
  sg13g2_a21oi_1 _18056_ (
    .A1(_02149_),
    .A2(_08360_),
    .B1(_08388_),
    .Y(_08361_)
  );
  sg13g2_a21oi_1 _18057_ (
    .A1(_00520_),
    .A2(_01267_),
    .B1(_03358_),
    .Y(_08362_)
  );
  sg13g2_nor2_1 _18058_ (
    .A(_08361_),
    .B(_08362_),
    .Y(_08363_)
  );
  sg13g2_o21ai_1 _18059_ (
    .A1(addr_i_3_),
    .A2(_08359_),
    .B1(_08363_),
    .Y(_08364_)
  );
  sg13g2_a21oi_1 _18060_ (
    .A1(_01273_),
    .A2(_00819_),
    .B1(addr_i_4_),
    .Y(_08366_)
  );
  sg13g2_a221oi_1 _18061_ (
    .A1(addr_i_3_),
    .A2(_00797_),
    .B1(_06129_),
    .B2(addr_i_2_),
    .C1(_08366_),
    .Y(_08367_)
  );
  sg13g2_nor2_1 _18062_ (
    .A(_01517_),
    .B(_08367_),
    .Y(_08368_)
  );
  sg13g2_o21ai_1 _18063_ (
    .A1(_03643_),
    .A2(_03742_),
    .B1(addr_i_4_),
    .Y(_08369_)
  );
  sg13g2_o21ai_1 _18064_ (
    .A1(_00226_),
    .A2(_04778_),
    .B1(_01674_),
    .Y(_08370_)
  );
  sg13g2_nand3_1 _18065_ (
    .A(_00618_),
    .B(_08369_),
    .C(_08370_),
    .Y(_08371_)
  );
  sg13g2_nor3_1 _18066_ (
    .A(addr_i_8_),
    .B(_08368_),
    .C(_08371_),
    .Y(_08372_)
  );
  sg13g2_a21oi_1 _18067_ (
    .A1(addr_i_8_),
    .A2(_08364_),
    .B1(_08372_),
    .Y(_08373_)
  );
  sg13g2_nor2_1 _18068_ (
    .A(_06939_),
    .B(_02069_),
    .Y(_08374_)
  );
  sg13g2_nand2_1 _18069_ (
    .A(_04904_),
    .B(_00679_),
    .Y(_08375_)
  );
  sg13g2_a22oi_1 _18070_ (
    .A1(addr_i_4_),
    .A2(_08375_),
    .B1(_00119_),
    .B2(addr_i_3_),
    .Y(_08378_)
  );
  sg13g2_a22oi_1 _18071_ (
    .A1(addr_i_3_),
    .A2(_08374_),
    .B1(_08378_),
    .B2(addr_i_2_),
    .Y(_08379_)
  );
  sg13g2_o21ai_1 _18072_ (
    .A1(_07348_),
    .A2(_09502_),
    .B1(addr_i_5_),
    .Y(_08380_)
  );
  sg13g2_o21ai_1 _18073_ (
    .A1(_01401_),
    .A2(_01567_),
    .B1(addr_i_3_),
    .Y(_08381_)
  );
  sg13g2_a21oi_1 _18074_ (
    .A1(_08380_),
    .A2(_08381_),
    .B1(_03281_),
    .Y(_08382_)
  );
  sg13g2_nor2_1 _18075_ (
    .A(_08379_),
    .B(_08382_),
    .Y(_08383_)
  );
  sg13g2_o21ai_1 _18076_ (
    .A1(_00056_),
    .A2(_03497_),
    .B1(_08383_),
    .Y(_08384_)
  );
  sg13g2_o21ai_1 _18077_ (
    .A1(_00297_),
    .A2(_03433_),
    .B1(addr_i_4_),
    .Y(_08385_)
  );
  sg13g2_and3_1 _18078_ (
    .A(_01008_),
    .B(_06439_),
    .C(_08385_),
    .X(_08386_)
  );
  sg13g2_o21ai_1 _18079_ (
    .A1(addr_i_3_),
    .A2(_00165_),
    .B1(_01120_),
    .Y(_08387_)
  );
  sg13g2_a21oi_1 _18080_ (
    .A1(_05596_),
    .A2(_08387_),
    .B1(_02777_),
    .Y(_08389_)
  );
  sg13g2_a22oi_1 _18081_ (
    .A1(_00645_),
    .A2(_05985_),
    .B1(_08389_),
    .B2(addr_i_2_),
    .Y(_08390_)
  );
  sg13g2_a22oi_1 _18082_ (
    .A1(addr_i_2_),
    .A2(_08386_),
    .B1(_08390_),
    .B2(addr_i_8_),
    .Y(_08391_)
  );
  sg13g2_a21oi_1 _18083_ (
    .A1(addr_i_8_),
    .A2(_08384_),
    .B1(_08391_),
    .Y(_08392_)
  );
  sg13g2_o21ai_1 _18084_ (
    .A1(addr_i_6_),
    .A2(_00759_),
    .B1(_00089_),
    .Y(_08393_)
  );
  sg13g2_a21oi_1 _18085_ (
    .A1(_04285_),
    .A2(_01152_),
    .B1(addr_i_3_),
    .Y(_08394_)
  );
  sg13g2_a22oi_1 _18086_ (
    .A1(addr_i_3_),
    .A2(_08393_),
    .B1(_08394_),
    .B2(_01837_),
    .Y(_08395_)
  );
  sg13g2_nor2_1 _18087_ (
    .A(_01095_),
    .B(_08395_),
    .Y(_08396_)
  );
  sg13g2_o21ai_1 _18088_ (
    .A1(_00965_),
    .A2(_00665_),
    .B1(_02150_),
    .Y(_08397_)
  );
  sg13g2_nand2_1 _18089_ (
    .A(addr_i_2_),
    .B(_08397_),
    .Y(_08398_)
  );
  sg13g2_nand3_1 _18090_ (
    .A(_01155_),
    .B(_00348_),
    .C(_01791_),
    .Y(_08400_)
  );
  sg13g2_nand3_1 _18091_ (
    .A(addr_i_8_),
    .B(_08398_),
    .C(_08400_),
    .Y(_08401_)
  );
  sg13g2_o21ai_1 _18092_ (
    .A1(_00946_),
    .A2(_07215_),
    .B1(addr_i_4_),
    .Y(_08402_)
  );
  sg13g2_a21oi_1 _18093_ (
    .A1(_01691_),
    .A2(_08402_),
    .B1(addr_i_5_),
    .Y(_08403_)
  );
  sg13g2_a21oi_1 _18094_ (
    .A1(_00687_),
    .A2(_01432_),
    .B1(_00965_),
    .Y(_08404_)
  );
  sg13g2_o21ai_1 _18095_ (
    .A1(_08403_),
    .A2(_08404_),
    .B1(addr_i_3_),
    .Y(_08405_)
  );
  sg13g2_a21oi_1 _18096_ (
    .A1(addr_i_5_),
    .A2(_00079_),
    .B1(_05025_),
    .Y(_08406_)
  );
  sg13g2_nor2_1 _18097_ (
    .A(_04528_),
    .B(_00099_),
    .Y(_08407_)
  );
  sg13g2_nor2_1 _18098_ (
    .A(_04384_),
    .B(_01264_),
    .Y(_08408_)
  );
  sg13g2_a22oi_1 _18099_ (
    .A1(addr_i_6_),
    .A2(_08407_),
    .B1(_08408_),
    .B2(addr_i_3_),
    .Y(_08409_)
  );
  sg13g2_o21ai_1 _18100_ (
    .A1(addr_i_6_),
    .A2(_08406_),
    .B1(_08409_),
    .Y(_08411_)
  );
  sg13g2_nand4_1 _18101_ (
    .A(_00629_),
    .B(_02082_),
    .C(_08405_),
    .D(_08411_),
    .Y(_08412_)
  );
  sg13g2_o21ai_1 _18102_ (
    .A1(_08396_),
    .A2(_08401_),
    .B1(_08412_),
    .Y(_08413_)
  );
  sg13g2_mux4_1 _18103_ (
    .A0(_08357_),
    .A1(_08373_),
    .A2(_08392_),
    .A3(_08413_),
    .S0(addr_i_9_),
    .S1(_03841_),
    .X(_08414_)
  );
  sg13g2_and2_1 _18104_ (
    .A(_00312_),
    .B(_08414_),
    .X(_08415_)
  );
  sg13g2_nor4_1 _18105_ (
    .A(_08179_),
    .B(_08252_),
    .C(_08331_),
    .D(_08415_),
    .Y(data_o_5_)
  );
  sg13g2_o21ai_1 _18106_ (
    .A1(_00087_),
    .A2(_02154_),
    .B1(addr_i_3_),
    .Y(_08416_)
  );
  sg13g2_nand2_1 _18107_ (
    .A(addr_i_5_),
    .B(_05769_),
    .Y(_08417_)
  );
  sg13g2_o21ai_1 _18108_ (
    .A1(_01508_),
    .A2(_07215_),
    .B1(_01653_),
    .Y(_08418_)
  );
  sg13g2_nand3_1 _18109_ (
    .A(_08416_),
    .B(_08417_),
    .C(_08418_),
    .Y(_08419_)
  );
  sg13g2_nand3_1 _18110_ (
    .A(addr_i_3_),
    .B(_00582_),
    .C(_01070_),
    .Y(_08421_)
  );
  sg13g2_a21oi_1 _18111_ (
    .A1(_01230_),
    .A2(_08421_),
    .B1(addr_i_6_),
    .Y(_08422_)
  );
  sg13g2_a22oi_1 _18112_ (
    .A1(_00191_),
    .A2(_08076_),
    .B1(_08422_),
    .B2(_03388_),
    .Y(_08423_)
  );
  sg13g2_a22oi_1 _18113_ (
    .A1(addr_i_4_),
    .A2(_08419_),
    .B1(_08423_),
    .B2(_06706_),
    .Y(_08424_)
  );
  sg13g2_a21o_1 _18114_ (
    .A1(_02471_),
    .A2(_07744_),
    .B1(addr_i_3_),
    .X(_08425_)
  );
  sg13g2_a21oi_1 _18115_ (
    .A1(_01203_),
    .A2(_08425_),
    .B1(_00146_),
    .Y(_08426_)
  );
  sg13g2_a22oi_1 _18116_ (
    .A1(_00239_),
    .A2(_01437_),
    .B1(_08426_),
    .B2(addr_i_6_),
    .Y(_08427_)
  );
  sg13g2_o21ai_1 _18117_ (
    .A1(addr_i_4_),
    .A2(_04238_),
    .B1(_08707_),
    .Y(_08428_)
  );
  sg13g2_a21oi_1 _18118_ (
    .A1(_00069_),
    .A2(_03783_),
    .B1(_00703_),
    .Y(_08429_)
  );
  sg13g2_a22oi_1 _18119_ (
    .A1(addr_i_2_),
    .A2(_08428_),
    .B1(_08429_),
    .B2(_00172_),
    .Y(_08430_)
  );
  sg13g2_a21oi_1 _18120_ (
    .A1(_01227_),
    .A2(_03572_),
    .B1(addr_i_8_),
    .Y(_08432_)
  );
  sg13g2_o21ai_1 _18121_ (
    .A1(_08427_),
    .A2(_08430_),
    .B1(_08432_),
    .Y(_08433_)
  );
  sg13g2_nand3b_1 _18122_ (
    .A_N(_08424_),
    .B(_05214_),
    .C(_08433_),
    .Y(_08434_)
  );
  sg13g2_o21ai_1 _18123_ (
    .A1(addr_i_2_),
    .A2(_01086_),
    .B1(_00200_),
    .Y(_08435_)
  );
  sg13g2_o21ai_1 _18124_ (
    .A1(addr_i_4_),
    .A2(_01094_),
    .B1(_08435_),
    .Y(_08436_)
  );
  sg13g2_o21ai_1 _18125_ (
    .A1(_02268_),
    .A2(_08436_),
    .B1(_00116_),
    .Y(_08437_)
  );
  sg13g2_nand2_1 _18126_ (
    .A(_02898_),
    .B(_03927_),
    .Y(_08438_)
  );
  sg13g2_a22oi_1 _18127_ (
    .A1(addr_i_3_),
    .A2(_08438_),
    .B1(_06276_),
    .B2(_00779_),
    .Y(_08439_)
  );
  sg13g2_a21oi_1 _18128_ (
    .A1(_01290_),
    .A2(_09476_),
    .B1(_00047_),
    .Y(_08440_)
  );
  sg13g2_a22oi_1 _18129_ (
    .A1(_00626_),
    .A2(_00727_),
    .B1(_01049_),
    .B2(_08440_),
    .Y(_08441_)
  );
  sg13g2_a221oi_1 _18130_ (
    .A1(_08437_),
    .A2(_08439_),
    .B1(_08441_),
    .B2(_05834_),
    .C1(_06706_),
    .Y(_08443_)
  );
  sg13g2_a21oi_1 _18131_ (
    .A1(_06088_),
    .A2(_01368_),
    .B1(_02472_),
    .Y(_08444_)
  );
  sg13g2_a21oi_1 _18132_ (
    .A1(_05402_),
    .A2(_06790_),
    .B1(_09348_),
    .Y(_08445_)
  );
  sg13g2_nor2_1 _18133_ (
    .A(addr_i_3_),
    .B(_08445_),
    .Y(_08446_)
  );
  sg13g2_a22oi_1 _18134_ (
    .A1(addr_i_3_),
    .A2(_02100_),
    .B1(_08444_),
    .B2(_08446_),
    .Y(_08447_)
  );
  sg13g2_and3_1 _18135_ (
    .A(_00870_),
    .B(_07359_),
    .C(_01843_),
    .X(_08448_)
  );
  sg13g2_a22oi_1 _18136_ (
    .A1(_00305_),
    .A2(_05873_),
    .B1(_08448_),
    .B2(addr_i_7_),
    .Y(_08449_)
  );
  sg13g2_a22oi_1 _18137_ (
    .A1(addr_i_7_),
    .A2(_08447_),
    .B1(_08449_),
    .B2(addr_i_8_),
    .Y(_08450_)
  );
  sg13g2_nand2b_1 _18138_ (
    .A_N(_08450_),
    .B(addr_i_9_),
    .Y(_08451_)
  );
  sg13g2_nor3_1 _18139_ (
    .A(_01499_),
    .B(_00031_),
    .C(_01246_),
    .Y(_08452_)
  );
  sg13g2_a22oi_1 _18140_ (
    .A1(_01892_),
    .A2(_04442_),
    .B1(_01612_),
    .B2(_08452_),
    .Y(_08454_)
  );
  sg13g2_o21ai_1 _18141_ (
    .A1(addr_i_3_),
    .A2(_00194_),
    .B1(_00077_),
    .Y(_08455_)
  );
  sg13g2_nand3_1 _18142_ (
    .A(addr_i_5_),
    .B(_01438_),
    .C(_02573_),
    .Y(_08456_)
  );
  sg13g2_o21ai_1 _18143_ (
    .A1(addr_i_5_),
    .A2(_08455_),
    .B1(_08456_),
    .Y(_08457_)
  );
  sg13g2_nand2_1 _18144_ (
    .A(addr_i_6_),
    .B(_00194_),
    .Y(_08458_)
  );
  sg13g2_o21ai_1 _18145_ (
    .A1(_02990_),
    .A2(_05737_),
    .B1(_08458_),
    .Y(_08459_)
  );
  sg13g2_nor2_1 _18146_ (
    .A(addr_i_6_),
    .B(_02418_),
    .Y(_08460_)
  );
  sg13g2_a22oi_1 _18147_ (
    .A1(_00497_),
    .A2(_08459_),
    .B1(_08460_),
    .B2(addr_i_2_),
    .Y(_08461_)
  );
  sg13g2_a21o_1 _18148_ (
    .A1(addr_i_2_),
    .A2(_08457_),
    .B1(_08461_),
    .X(_08462_)
  );
  sg13g2_o21ai_1 _18149_ (
    .A1(_04439_),
    .A2(_00057_),
    .B1(_00060_),
    .Y(_08463_)
  );
  sg13g2_o21ai_1 _18150_ (
    .A1(_00899_),
    .A2(_02744_),
    .B1(_08463_),
    .Y(_08465_)
  );
  sg13g2_o21ai_1 _18151_ (
    .A1(_00305_),
    .A2(_00057_),
    .B1(addr_i_5_),
    .Y(_08466_)
  );
  sg13g2_nand3_1 _18152_ (
    .A(addr_i_4_),
    .B(addr_i_6_),
    .C(_02577_),
    .Y(_08467_)
  );
  sg13g2_a21oi_1 _18153_ (
    .A1(_08466_),
    .A2(_08467_),
    .B1(_00315_),
    .Y(_08468_)
  );
  sg13g2_a22oi_1 _18154_ (
    .A1(_00068_),
    .A2(_08465_),
    .B1(_08468_),
    .B2(_02368_),
    .Y(_08469_)
  );
  sg13g2_a22oi_1 _18155_ (
    .A1(_08454_),
    .A2(_08462_),
    .B1(addr_i_10_),
    .B2(_08469_),
    .Y(_08470_)
  );
  sg13g2_o21ai_1 _18156_ (
    .A1(_08443_),
    .A2(_08451_),
    .B1(_08470_),
    .Y(_08471_)
  );
  sg13g2_nand2_1 _18157_ (
    .A(addr_i_3_),
    .B(_05960_),
    .Y(_08472_)
  );
  sg13g2_a21oi_1 _18158_ (
    .A1(_03944_),
    .A2(_08472_),
    .B1(_01279_),
    .Y(_08473_)
  );
  sg13g2_a21oi_1 _18159_ (
    .A1(_01227_),
    .A2(_03262_),
    .B1(_08473_),
    .Y(_08474_)
  );
  sg13g2_a22oi_1 _18160_ (
    .A1(_00159_),
    .A2(_00820_),
    .B1(_02265_),
    .B2(_00588_),
    .Y(_08476_)
  );
  sg13g2_o21ai_1 _18161_ (
    .A1(_00569_),
    .A2(_03936_),
    .B1(_08476_),
    .Y(_08477_)
  );
  sg13g2_o21ai_1 _18162_ (
    .A1(_01391_),
    .A2(_08474_),
    .B1(_08477_),
    .Y(_08478_)
  );
  sg13g2_a22oi_1 _18163_ (
    .A1(_01277_),
    .A2(_01437_),
    .B1(_05645_),
    .B2(_00083_),
    .Y(_08479_)
  );
  sg13g2_a22oi_1 _18164_ (
    .A1(_00827_),
    .A2(_09486_),
    .B1(_00959_),
    .B2(addr_i_4_),
    .Y(_08480_)
  );
  sg13g2_o21ai_1 _18165_ (
    .A1(_08479_),
    .A2(_08480_),
    .B1(_02349_),
    .Y(_08481_)
  );
  sg13g2_a21oi_1 _18166_ (
    .A1(_00930_),
    .A2(_00926_),
    .B1(addr_i_5_),
    .Y(_08482_)
  );
  sg13g2_a21oi_1 _18167_ (
    .A1(_00930_),
    .A2(_01834_),
    .B1(addr_i_3_),
    .Y(_08483_)
  );
  sg13g2_o21ai_1 _18168_ (
    .A1(_08482_),
    .A2(_08483_),
    .B1(_02796_),
    .Y(_08484_)
  );
  sg13g2_o21ai_1 _18169_ (
    .A1(_02578_),
    .A2(_00764_),
    .B1(_08484_),
    .Y(_08485_)
  );
  sg13g2_a21oi_1 _18170_ (
    .A1(addr_i_3_),
    .A2(_08481_),
    .B1(_08485_),
    .Y(_08488_)
  );
  sg13g2_nor2_1 _18171_ (
    .A(addr_i_8_),
    .B(_08488_),
    .Y(_08489_)
  );
  sg13g2_o21ai_1 _18172_ (
    .A1(_08478_),
    .A2(_08489_),
    .B1(_01176_),
    .Y(_08490_)
  );
  sg13g2_nand4_1 _18173_ (
    .A(addr_i_11_),
    .B(_08434_),
    .C(_08471_),
    .D(_08490_),
    .Y(_08491_)
  );
  sg13g2_nand2_1 _18174_ (
    .A(_00505_),
    .B(_09494_),
    .Y(_08492_)
  );
  sg13g2_nand2_1 _18175_ (
    .A(_00105_),
    .B(_08492_),
    .Y(_08493_)
  );
  sg13g2_o21ai_1 _18176_ (
    .A1(addr_i_2_),
    .A2(_03336_),
    .B1(_09260_),
    .Y(_08494_)
  );
  sg13g2_a221oi_1 _18177_ (
    .A1(addr_i_2_),
    .A2(_08493_),
    .B1(_08494_),
    .B2(addr_i_7_),
    .C1(_04281_),
    .Y(_08495_)
  );
  sg13g2_a22oi_1 _18178_ (
    .A1(addr_i_4_),
    .A2(_03112_),
    .B1(_01380_),
    .B2(_01837_),
    .Y(_08496_)
  );
  sg13g2_a221oi_1 _18179_ (
    .A1(_03142_),
    .A2(_06372_),
    .B1(_08496_),
    .B2(addr_i_7_),
    .C1(addr_i_3_),
    .Y(_08497_)
  );
  sg13g2_a21oi_1 _18180_ (
    .A1(_01365_),
    .A2(_00301_),
    .B1(_08497_),
    .Y(_08499_)
  );
  sg13g2_o21ai_1 _18181_ (
    .A1(_00048_),
    .A2(_08495_),
    .B1(_08499_),
    .Y(_08500_)
  );
  sg13g2_a21oi_1 _18182_ (
    .A1(_01350_),
    .A2(_08500_),
    .B1(addr_i_11_),
    .Y(_08501_)
  );
  sg13g2_nand2_1 _18183_ (
    .A(_01616_),
    .B(_00645_),
    .Y(_08502_)
  );
  sg13g2_o21ai_1 _18184_ (
    .A1(_00051_),
    .A2(_00315_),
    .B1(_08502_),
    .Y(_08503_)
  );
  sg13g2_nand3_1 _18185_ (
    .A(_00091_),
    .B(_00716_),
    .C(_03660_),
    .Y(_08504_)
  );
  sg13g2_nand3_1 _18186_ (
    .A(addr_i_6_),
    .B(_00522_),
    .C(_02840_),
    .Y(_08505_)
  );
  sg13g2_nand3_1 _18187_ (
    .A(addr_i_7_),
    .B(_08504_),
    .C(_08505_),
    .Y(_08506_)
  );
  sg13g2_a21oi_1 _18188_ (
    .A1(_00656_),
    .A2(_08506_),
    .B1(addr_i_2_),
    .Y(_08507_)
  );
  sg13g2_a21o_1 _18189_ (
    .A1(addr_i_4_),
    .A2(_08503_),
    .B1(_08507_),
    .X(_08508_)
  );
  sg13g2_nor3_1 _18190_ (
    .A(addr_i_2_),
    .B(_01815_),
    .C(_02781_),
    .Y(_08510_)
  );
  sg13g2_nand2_1 _18191_ (
    .A(_00064_),
    .B(_01920_),
    .Y(_08511_)
  );
  sg13g2_a21oi_1 _18192_ (
    .A1(_03575_),
    .A2(_08511_),
    .B1(_01095_),
    .Y(_08512_)
  );
  sg13g2_o21ai_1 _18193_ (
    .A1(_08510_),
    .A2(_08512_),
    .B1(addr_i_3_),
    .Y(_08513_)
  );
  sg13g2_o21ai_1 _18194_ (
    .A1(_00827_),
    .A2(_06198_),
    .B1(addr_i_4_),
    .Y(_08514_)
  );
  sg13g2_nor3_1 _18195_ (
    .A(_00015_),
    .B(_01514_),
    .C(_05112_),
    .Y(_08515_)
  );
  sg13g2_o21ai_1 _18196_ (
    .A1(addr_i_4_),
    .A2(_03465_),
    .B1(_07625_),
    .Y(_08516_)
  );
  sg13g2_o21ai_1 _18197_ (
    .A1(addr_i_8_),
    .A2(_01265_),
    .B1(addr_i_7_),
    .Y(_08517_)
  );
  sg13g2_a221oi_1 _18198_ (
    .A1(_08514_),
    .A2(_08515_),
    .B1(_08516_),
    .B2(_01519_),
    .C1(_08517_),
    .Y(_08518_)
  );
  sg13g2_a21oi_1 _18199_ (
    .A1(_00566_),
    .A2(_00470_),
    .B1(addr_i_8_),
    .Y(_08519_)
  );
  sg13g2_a21oi_1 _18200_ (
    .A1(_08930_),
    .A2(_02781_),
    .B1(addr_i_3_),
    .Y(_08521_)
  );
  sg13g2_o21ai_1 _18201_ (
    .A1(_08519_),
    .A2(_08521_),
    .B1(_09271_),
    .Y(_08522_)
  );
  sg13g2_a21oi_1 _18202_ (
    .A1(_01019_),
    .A2(_06408_),
    .B1(_00067_),
    .Y(_08523_)
  );
  sg13g2_o21ai_1 _18203_ (
    .A1(addr_i_3_),
    .A2(_02388_),
    .B1(_03226_),
    .Y(_08524_)
  );
  sg13g2_a21oi_1 _18204_ (
    .A1(addr_i_8_),
    .A2(_00550_),
    .B1(_06441_),
    .Y(_08525_)
  );
  sg13g2_o21ai_1 _18205_ (
    .A1(_08951_),
    .A2(_08525_),
    .B1(_06406_),
    .Y(_08526_)
  );
  sg13g2_a22oi_1 _18206_ (
    .A1(addr_i_8_),
    .A2(_08524_),
    .B1(_08526_),
    .B2(addr_i_2_),
    .Y(_08527_)
  );
  sg13g2_a21oi_1 _18207_ (
    .A1(_08522_),
    .A2(_08523_),
    .B1(_08527_),
    .Y(_08528_)
  );
  sg13g2_a22oi_1 _18208_ (
    .A1(_07547_),
    .A2(_06405_),
    .B1(_08528_),
    .B2(addr_i_7_),
    .Y(_08529_)
  );
  sg13g2_a22oi_1 _18209_ (
    .A1(_08513_),
    .A2(_08518_),
    .B1(_02221_),
    .B2(_08529_),
    .Y(_08530_)
  );
  sg13g2_nand2_1 _18210_ (
    .A(_02887_),
    .B(_01087_),
    .Y(_08532_)
  );
  sg13g2_o21ai_1 _18211_ (
    .A1(addr_i_2_),
    .A2(_07237_),
    .B1(addr_i_3_),
    .Y(_08533_)
  );
  sg13g2_a21oi_1 _18212_ (
    .A1(_01912_),
    .A2(_08533_),
    .B1(addr_i_6_),
    .Y(_08534_)
  );
  sg13g2_a22oi_1 _18213_ (
    .A1(_00115_),
    .A2(_08532_),
    .B1(_08534_),
    .B2(_06276_),
    .Y(_08535_)
  );
  sg13g2_a21oi_1 _18214_ (
    .A1(_04528_),
    .A2(_00676_),
    .B1(_03632_),
    .Y(_08536_)
  );
  sg13g2_a21o_1 _18215_ (
    .A1(_01636_),
    .A2(_00785_),
    .B1(_00711_),
    .X(_08537_)
  );
  sg13g2_o21ai_1 _18216_ (
    .A1(addr_i_3_),
    .A2(_08536_),
    .B1(_08537_),
    .Y(_08538_)
  );
  sg13g2_a21oi_1 _18217_ (
    .A1(_00368_),
    .A2(_03258_),
    .B1(_02076_),
    .Y(_08539_)
  );
  sg13g2_a21oi_1 _18218_ (
    .A1(addr_i_7_),
    .A2(_08538_),
    .B1(_08539_),
    .Y(_08540_)
  );
  sg13g2_o21ai_1 _18219_ (
    .A1(addr_i_7_),
    .A2(_08535_),
    .B1(_08540_),
    .Y(_08541_)
  );
  sg13g2_a22oi_1 _18220_ (
    .A1(addr_i_3_),
    .A2(_06790_),
    .B1(_00746_),
    .B2(_00743_),
    .Y(_08543_)
  );
  sg13g2_nor3_1 _18221_ (
    .A(addr_i_4_),
    .B(_06497_),
    .C(_00857_),
    .Y(_08544_)
  );
  sg13g2_a22oi_1 _18222_ (
    .A1(addr_i_4_),
    .A2(_08543_),
    .B1(_08544_),
    .B2(_07403_),
    .Y(_08545_)
  );
  sg13g2_nor2_1 _18223_ (
    .A(_00011_),
    .B(_03245_),
    .Y(_08546_)
  );
  sg13g2_a22oi_1 _18224_ (
    .A1(addr_i_3_),
    .A2(_08546_),
    .B1(_02057_),
    .B2(_03652_),
    .Y(_08547_)
  );
  sg13g2_o21ai_1 _18225_ (
    .A1(addr_i_4_),
    .A2(_03979_),
    .B1(_01666_),
    .Y(_08548_)
  );
  sg13g2_o21ai_1 _18226_ (
    .A1(_08547_),
    .A2(_08548_),
    .B1(addr_i_9_),
    .Y(_08549_)
  );
  sg13g2_a22oi_1 _18227_ (
    .A1(_00367_),
    .A2(_08541_),
    .B1(_08545_),
    .B2(_08549_),
    .Y(_08550_)
  );
  sg13g2_nand2_1 _18228_ (
    .A(_00840_),
    .B(_07087_),
    .Y(_08551_)
  );
  sg13g2_nand3_1 _18229_ (
    .A(addr_i_3_),
    .B(_03325_),
    .C(_04077_),
    .Y(_08552_)
  );
  sg13g2_a21oi_1 _18230_ (
    .A1(_01397_),
    .A2(_08552_),
    .B1(_03919_),
    .Y(_08554_)
  );
  sg13g2_a22oi_1 _18231_ (
    .A1(_03993_),
    .A2(_03772_),
    .B1(_08554_),
    .B2(_05218_),
    .Y(_08555_)
  );
  sg13g2_a22oi_1 _18232_ (
    .A1(_01788_),
    .A2(_08551_),
    .B1(_08555_),
    .B2(_03617_),
    .Y(_08556_)
  );
  sg13g2_nand2_1 _18233_ (
    .A(_00479_),
    .B(_01754_),
    .Y(_08557_)
  );
  sg13g2_nand2_1 _18234_ (
    .A(_01436_),
    .B(_08453_),
    .Y(_08558_)
  );
  sg13g2_a21o_1 _18235_ (
    .A1(_08557_),
    .A2(_08558_),
    .B1(_00200_),
    .X(_08559_)
  );
  sg13g2_a21oi_1 _18236_ (
    .A1(_00314_),
    .A2(_08559_),
    .B1(_08830_),
    .Y(_08560_)
  );
  sg13g2_o21ai_1 _18237_ (
    .A1(_05568_),
    .A2(_00415_),
    .B1(_00616_),
    .Y(_08561_)
  );
  sg13g2_a21oi_1 _18238_ (
    .A1(_03564_),
    .A2(_08561_),
    .B1(_07614_),
    .Y(_08562_)
  );
  sg13g2_nor4_1 _18239_ (
    .A(addr_i_9_),
    .B(_08556_),
    .C(_08560_),
    .D(_08562_),
    .Y(_08563_)
  );
  sg13g2_nor3_1 _18240_ (
    .A(addr_i_10_),
    .B(_08550_),
    .C(_08563_),
    .Y(_08565_)
  );
  sg13g2_a22oi_1 _18241_ (
    .A1(_01613_),
    .A2(_08508_),
    .B1(_08530_),
    .B2(_08565_),
    .Y(_08566_)
  );
  sg13g2_a21oi_1 _18242_ (
    .A1(_08501_),
    .A2(_08566_),
    .B1(addr_i_12_),
    .Y(_08567_)
  );
  sg13g2_a21o_1 _18243_ (
    .A1(addr_i_4_),
    .A2(_00275_),
    .B1(_03914_),
    .X(_08568_)
  );
  sg13g2_a21oi_1 _18244_ (
    .A1(_01367_),
    .A2(_01230_),
    .B1(addr_i_4_),
    .Y(_08569_)
  );
  sg13g2_a221oi_1 _18245_ (
    .A1(_01747_),
    .A2(_00745_),
    .B1(_08568_),
    .B2(addr_i_3_),
    .C1(_08569_),
    .Y(_08570_)
  );
  sg13g2_nor3_1 _18246_ (
    .A(addr_i_4_),
    .B(_03245_),
    .C(_02514_),
    .Y(_08571_)
  );
  sg13g2_a21oi_1 _18247_ (
    .A1(_07370_),
    .A2(_07736_),
    .B1(_08571_),
    .Y(_08572_)
  );
  sg13g2_a21oi_1 _18248_ (
    .A1(_02694_),
    .A2(_02898_),
    .B1(addr_i_3_),
    .Y(_08573_)
  );
  sg13g2_o21ai_1 _18249_ (
    .A1(_08572_),
    .A2(_08573_),
    .B1(addr_i_7_),
    .Y(_08574_)
  );
  sg13g2_nand2_1 _18250_ (
    .A(_08570_),
    .B(_08574_),
    .Y(_08576_)
  );
  sg13g2_a21oi_1 _18251_ (
    .A1(addr_i_3_),
    .A2(_08407_),
    .B1(_08598_),
    .Y(_08577_)
  );
  sg13g2_o21ai_1 _18252_ (
    .A1(addr_i_6_),
    .A2(_08577_),
    .B1(_06735_),
    .Y(_08578_)
  );
  sg13g2_a21oi_1 _18253_ (
    .A1(addr_i_3_),
    .A2(_04355_),
    .B1(_01380_),
    .Y(_08579_)
  );
  sg13g2_nor4_1 _18254_ (
    .A(addr_i_3_),
    .B(_08653_),
    .C(_00032_),
    .D(_04539_),
    .Y(_08580_)
  );
  sg13g2_a22oi_1 _18255_ (
    .A1(_01567_),
    .A2(_04713_),
    .B1(_08580_),
    .B2(_01611_),
    .Y(_08581_)
  );
  sg13g2_o21ai_1 _18256_ (
    .A1(_00324_),
    .A2(_08579_),
    .B1(_08581_),
    .Y(_08582_)
  );
  sg13g2_nor2_1 _18257_ (
    .A(_00051_),
    .B(_01831_),
    .Y(_08583_)
  );
  sg13g2_a22oi_1 _18258_ (
    .A1(_01324_),
    .A2(_08578_),
    .B1(_08582_),
    .B2(_08583_),
    .Y(_08584_)
  );
  sg13g2_a22oi_1 _18259_ (
    .A1(_00423_),
    .A2(_08576_),
    .B1(_08584_),
    .B2(_03841_),
    .Y(_08585_)
  );
  sg13g2_o21ai_1 _18260_ (
    .A1(_00386_),
    .A2(_00234_),
    .B1(_01500_),
    .Y(_08587_)
  );
  sg13g2_a21oi_1 _18261_ (
    .A1(addr_i_6_),
    .A2(_04494_),
    .B1(_02387_),
    .Y(_08588_)
  );
  sg13g2_o21ai_1 _18262_ (
    .A1(_02428_),
    .A2(_08588_),
    .B1(addr_i_2_),
    .Y(_08589_)
  );
  sg13g2_a21oi_1 _18263_ (
    .A1(_08587_),
    .A2(_08589_),
    .B1(_01279_),
    .Y(_08590_)
  );
  sg13g2_o21ai_1 _18264_ (
    .A1(_01086_),
    .A2(_08299_),
    .B1(addr_i_3_),
    .Y(_08591_)
  );
  sg13g2_a21oi_1 _18265_ (
    .A1(_01267_),
    .A2(_08591_),
    .B1(_01475_),
    .Y(_08592_)
  );
  sg13g2_a22oi_1 _18266_ (
    .A1(_00500_),
    .A2(_03572_),
    .B1(_08590_),
    .B2(_08592_),
    .Y(_08593_)
  );
  sg13g2_a21oi_1 _18267_ (
    .A1(_08874_),
    .A2(_03445_),
    .B1(_01663_),
    .Y(_08594_)
  );
  sg13g2_a221oi_1 _18268_ (
    .A1(_09050_),
    .A2(_07492_),
    .B1(_00571_),
    .B2(_02369_),
    .C1(_08696_),
    .Y(_08595_)
  );
  sg13g2_a22oi_1 _18269_ (
    .A1(_04284_),
    .A2(_08111_),
    .B1(_08122_),
    .B2(addr_i_5_),
    .Y(_08596_)
  );
  sg13g2_nor2_1 _18270_ (
    .A(_08595_),
    .B(_08596_),
    .Y(_08599_)
  );
  sg13g2_a21oi_1 _18271_ (
    .A1(_09486_),
    .A2(_00157_),
    .B1(_08599_),
    .Y(_08600_)
  );
  sg13g2_o21ai_1 _18272_ (
    .A1(addr_i_3_),
    .A2(_01228_),
    .B1(_00333_),
    .Y(_08601_)
  );
  sg13g2_a22oi_1 _18273_ (
    .A1(addr_i_4_),
    .A2(_08601_),
    .B1(_00898_),
    .B2(addr_i_2_),
    .Y(_08602_)
  );
  sg13g2_a22oi_1 _18274_ (
    .A1(addr_i_2_),
    .A2(_08600_),
    .B1(_08602_),
    .B2(_00113_),
    .Y(_08603_)
  );
  sg13g2_nor3_1 _18275_ (
    .A(_04705_),
    .B(_08594_),
    .C(_08603_),
    .Y(_08604_)
  );
  sg13g2_o21ai_1 _18276_ (
    .A1(addr_i_8_),
    .A2(_08593_),
    .B1(_08604_),
    .Y(_08605_)
  );
  sg13g2_o21ai_1 _18277_ (
    .A1(_03980_),
    .A2(_01031_),
    .B1(_03348_),
    .Y(_08606_)
  );
  sg13g2_o21ai_1 _18278_ (
    .A1(_07879_),
    .A2(_02490_),
    .B1(_01277_),
    .Y(_08607_)
  );
  sg13g2_nand3b_1 _18279_ (
    .A_N(_04681_),
    .B(_08606_),
    .C(_08607_),
    .Y(_08608_)
  );
  sg13g2_o21ai_1 _18280_ (
    .A1(_00616_),
    .A2(_00127_),
    .B1(addr_i_5_),
    .Y(_08610_)
  );
  sg13g2_a21oi_1 _18281_ (
    .A1(_02467_),
    .A2(_08610_),
    .B1(_01099_),
    .Y(_08611_)
  );
  sg13g2_a22oi_1 _18282_ (
    .A1(_00708_),
    .A2(_08608_),
    .B1(_08611_),
    .B2(addr_i_9_),
    .Y(_08612_)
  );
  sg13g2_a21oi_1 _18283_ (
    .A1(addr_i_4_),
    .A2(_03262_),
    .B1(_05306_),
    .Y(_08613_)
  );
  sg13g2_o21ai_1 _18284_ (
    .A1(addr_i_3_),
    .A2(_08613_),
    .B1(_07877_),
    .Y(_08614_)
  );
  sg13g2_o21ai_1 _18285_ (
    .A1(_08475_),
    .A2(_07601_),
    .B1(_00083_),
    .Y(_08615_)
  );
  sg13g2_a21o_1 _18286_ (
    .A1(_09415_),
    .A2(_02285_),
    .B1(_04461_),
    .X(_08616_)
  );
  sg13g2_a21oi_1 _18287_ (
    .A1(_08615_),
    .A2(_08616_),
    .B1(_00600_),
    .Y(_08617_)
  );
  sg13g2_a21oi_1 _18288_ (
    .A1(_01861_),
    .A2(_08614_),
    .B1(_08617_),
    .Y(_08618_)
  );
  sg13g2_a21oi_1 _18289_ (
    .A1(_00549_),
    .A2(_02920_),
    .B1(addr_i_3_),
    .Y(_08619_)
  );
  sg13g2_a21oi_1 _18290_ (
    .A1(addr_i_3_),
    .A2(_01998_),
    .B1(_08619_),
    .Y(_08621_)
  );
  sg13g2_a21oi_1 _18291_ (
    .A1(_01420_),
    .A2(_04367_),
    .B1(_04837_),
    .Y(_08622_)
  );
  sg13g2_o21ai_1 _18292_ (
    .A1(addr_i_5_),
    .A2(_08621_),
    .B1(_08622_),
    .Y(_08623_)
  );
  sg13g2_a21oi_1 _18293_ (
    .A1(addr_i_6_),
    .A2(_00582_),
    .B1(addr_i_4_),
    .Y(_08624_)
  );
  sg13g2_o21ai_1 _18294_ (
    .A1(addr_i_5_),
    .A2(_01439_),
    .B1(_00244_),
    .Y(_08625_)
  );
  sg13g2_o21ai_1 _18295_ (
    .A1(_08166_),
    .A2(_03245_),
    .B1(addr_i_3_),
    .Y(_08626_)
  );
  sg13g2_nand2_1 _18296_ (
    .A(_08625_),
    .B(_08626_),
    .Y(_08627_)
  );
  sg13g2_a21oi_1 _18297_ (
    .A1(_01160_),
    .A2(_02683_),
    .B1(_08266_),
    .Y(_08628_)
  );
  sg13g2_nor4_1 _18298_ (
    .A(_00860_),
    .B(_08624_),
    .C(_08627_),
    .D(_08628_),
    .Y(_08629_)
  );
  sg13g2_a22oi_1 _18299_ (
    .A1(_00708_),
    .A2(_08623_),
    .B1(_08629_),
    .B2(_04705_),
    .Y(_08630_)
  );
  sg13g2_a21oi_1 _18300_ (
    .A1(_00616_),
    .A2(_00770_),
    .B1(_03648_),
    .Y(_08632_)
  );
  sg13g2_a22oi_1 _18301_ (
    .A1(addr_i_3_),
    .A2(_03942_),
    .B1(_03720_),
    .B2(_02441_),
    .Y(_08633_)
  );
  sg13g2_mux2_1 _18302_ (
    .A0(_08632_),
    .A1(_08633_),
    .S(addr_i_5_),
    .X(_08634_)
  );
  sg13g2_nand3_1 _18303_ (
    .A(addr_i_8_),
    .B(_00852_),
    .C(_08634_),
    .Y(_08635_)
  );
  sg13g2_a22oi_1 _18304_ (
    .A1(_01450_),
    .A2(_01179_),
    .B1(_02228_),
    .B2(_01114_),
    .Y(_08636_)
  );
  sg13g2_a221oi_1 _18305_ (
    .A1(_00990_),
    .A2(_02107_),
    .B1(_03170_),
    .B2(_01970_),
    .C1(addr_i_4_),
    .Y(_08637_)
  );
  sg13g2_o21ai_1 _18306_ (
    .A1(_08636_),
    .A2(_08637_),
    .B1(_03617_),
    .Y(_08638_)
  );
  sg13g2_nand3_1 _18307_ (
    .A(addr_i_7_),
    .B(_08635_),
    .C(_08638_),
    .Y(_08639_)
  );
  sg13g2_a221oi_1 _18308_ (
    .A1(_08612_),
    .A2(_08618_),
    .B1(_08630_),
    .B2(_08639_),
    .C1(addr_i_10_),
    .Y(_08640_)
  );
  sg13g2_a21oi_1 _18309_ (
    .A1(_08585_),
    .A2(_08605_),
    .B1(_08640_),
    .Y(_08641_)
  );
  sg13g2_o21ai_1 _18310_ (
    .A1(_00204_),
    .A2(_00206_),
    .B1(_00068_),
    .Y(_08643_)
  );
  sg13g2_nand2_1 _18311_ (
    .A(_07288_),
    .B(_08643_),
    .Y(_08644_)
  );
  sg13g2_nor2_1 _18312_ (
    .A(_09315_),
    .B(_02672_),
    .Y(_08645_)
  );
  sg13g2_nand2_1 _18313_ (
    .A(_00852_),
    .B(_04145_),
    .Y(_08646_)
  );
  sg13g2_nor2_1 _18314_ (
    .A(_01007_),
    .B(_02505_),
    .Y(_08647_)
  );
  sg13g2_a22oi_1 _18315_ (
    .A1(_04251_),
    .A2(_08646_),
    .B1(_08647_),
    .B2(addr_i_7_),
    .Y(_08648_)
  );
  sg13g2_a22oi_1 _18316_ (
    .A1(addr_i_7_),
    .A2(_01656_),
    .B1(_08648_),
    .B2(addr_i_9_),
    .Y(_08649_)
  );
  sg13g2_o21ai_1 _18317_ (
    .A1(_08645_),
    .A2(_08649_),
    .B1(addr_i_8_),
    .Y(_08650_)
  );
  sg13g2_nor2_1 _18318_ (
    .A(_09513_),
    .B(_00405_),
    .Y(_08651_)
  );
  sg13g2_a21oi_1 _18319_ (
    .A1(addr_i_3_),
    .A2(_07969_),
    .B1(_08651_),
    .Y(_08652_)
  );
  sg13g2_o21ai_1 _18320_ (
    .A1(_01276_),
    .A2(_06541_),
    .B1(_01120_),
    .Y(_08654_)
  );
  sg13g2_a21oi_1 _18321_ (
    .A1(_02187_),
    .A2(_08654_),
    .B1(addr_i_3_),
    .Y(_08655_)
  );
  sg13g2_o21ai_1 _18322_ (
    .A1(_08475_),
    .A2(_08655_),
    .B1(addr_i_7_),
    .Y(_08656_)
  );
  sg13g2_o21ai_1 _18323_ (
    .A1(addr_i_2_),
    .A2(_08652_),
    .B1(_08656_),
    .Y(_08657_)
  );
  sg13g2_nand3_1 _18324_ (
    .A(addr_i_7_),
    .B(_03465_),
    .C(_08774_),
    .Y(_08658_)
  );
  sg13g2_nand2_1 _18325_ (
    .A(_01615_),
    .B(_01656_),
    .Y(_08659_)
  );
  sg13g2_a21oi_1 _18326_ (
    .A1(_08658_),
    .A2(_08659_),
    .B1(_09315_),
    .Y(_08660_)
  );
  sg13g2_a21oi_1 _18327_ (
    .A1(_00423_),
    .A2(_08657_),
    .B1(_08660_),
    .Y(_08661_)
  );
  sg13g2_a21oi_1 _18328_ (
    .A1(_08650_),
    .A2(_08661_),
    .B1(addr_i_10_),
    .Y(_08662_)
  );
  sg13g2_a22oi_1 _18329_ (
    .A1(_03084_),
    .A2(_08644_),
    .B1(_08662_),
    .B2(_07319_),
    .Y(_08663_)
  );
  sg13g2_a22oi_1 _18330_ (
    .A1(_03051_),
    .A2(_08641_),
    .B1(_08663_),
    .B2(_00812_),
    .Y(_08665_)
  );
  sg13g2_a21o_1 _18331_ (
    .A1(_08491_),
    .A2(_08567_),
    .B1(_08665_),
    .X(data_o_6_)
  );
  sg13g2_nand2_1 _18332_ (
    .A(_00316_),
    .B(_08852_),
    .Y(_08666_)
  );
  sg13g2_nand3_1 _18333_ (
    .A(_07284_),
    .B(_02546_),
    .C(_08666_),
    .Y(_08667_)
  );
  sg13g2_a21oi_1 _18334_ (
    .A1(addr_i_3_),
    .A2(_08796_),
    .B1(_06099_),
    .Y(_08668_)
  );
  sg13g2_nor2_1 _18335_ (
    .A(_01603_),
    .B(_08668_),
    .Y(_08669_)
  );
  sg13g2_a21oi_1 _18336_ (
    .A1(addr_i_5_),
    .A2(_08667_),
    .B1(_08669_),
    .Y(_08670_)
  );
  sg13g2_nor2_1 _18337_ (
    .A(_01276_),
    .B(_01048_),
    .Y(_08671_)
  );
  sg13g2_o21ai_1 _18338_ (
    .A1(addr_i_3_),
    .A2(_08671_),
    .B1(_01224_),
    .Y(_08672_)
  );
  sg13g2_nand2_1 _18339_ (
    .A(_04108_),
    .B(_01164_),
    .Y(_08673_)
  );
  sg13g2_a21oi_1 _18340_ (
    .A1(_08232_),
    .A2(_08673_),
    .B1(_00115_),
    .Y(_08675_)
  );
  sg13g2_o21ai_1 _18341_ (
    .A1(_00930_),
    .A2(_07769_),
    .B1(_06684_),
    .Y(_08676_)
  );
  sg13g2_a22oi_1 _18342_ (
    .A1(_01517_),
    .A2(_08672_),
    .B1(_08675_),
    .B2(_08676_),
    .Y(_08677_)
  );
  sg13g2_o21ai_1 _18343_ (
    .A1(_08399_),
    .A2(_08670_),
    .B1(_08677_),
    .Y(_08678_)
  );
  sg13g2_a21oi_1 _18344_ (
    .A1(_02815_),
    .A2(_01912_),
    .B1(addr_i_3_),
    .Y(_08679_)
  );
  sg13g2_a22oi_1 _18345_ (
    .A1(addr_i_4_),
    .A2(_07025_),
    .B1(_09094_),
    .B2(_08679_),
    .Y(_08680_)
  );
  sg13g2_nor2_1 _18346_ (
    .A(_08785_),
    .B(_02808_),
    .Y(_08681_)
  );
  sg13g2_o21ai_1 _18347_ (
    .A1(_07248_),
    .A2(_08681_),
    .B1(_03281_),
    .Y(_08682_)
  );
  sg13g2_nor3_1 _18348_ (
    .A(_04307_),
    .B(_00319_),
    .C(_02312_),
    .Y(_08683_)
  );
  sg13g2_a21oi_1 _18349_ (
    .A1(_08682_),
    .A2(_08683_),
    .B1(_01559_),
    .Y(_08684_)
  );
  sg13g2_o21ai_1 _18350_ (
    .A1(_06905_),
    .A2(_08680_),
    .B1(_08684_),
    .Y(_08686_)
  );
  sg13g2_o21ai_1 _18351_ (
    .A1(_02744_),
    .A2(_02528_),
    .B1(_01118_),
    .Y(_08687_)
  );
  sg13g2_a22oi_1 _18352_ (
    .A1(addr_i_6_),
    .A2(_05557_),
    .B1(_02954_),
    .B2(_08687_),
    .Y(_08688_)
  );
  sg13g2_a21o_1 _18353_ (
    .A1(_08678_),
    .A2(_08686_),
    .B1(_08688_),
    .X(_08689_)
  );
  sg13g2_a21oi_1 _18354_ (
    .A1(addr_i_7_),
    .A2(_03061_),
    .B1(_01837_),
    .Y(_08690_)
  );
  sg13g2_a21oi_1 _18355_ (
    .A1(_00516_),
    .A2(_04715_),
    .B1(_00648_),
    .Y(_08691_)
  );
  sg13g2_a21oi_1 _18356_ (
    .A1(_00261_),
    .A2(_06983_),
    .B1(_08691_),
    .Y(_08692_)
  );
  sg13g2_a21oi_1 _18357_ (
    .A1(_08690_),
    .A2(_08692_),
    .B1(addr_i_3_),
    .Y(_08693_)
  );
  sg13g2_nand2_1 _18358_ (
    .A(_00006_),
    .B(_01570_),
    .Y(_08694_)
  );
  sg13g2_a22oi_1 _18359_ (
    .A1(addr_i_4_),
    .A2(_02426_),
    .B1(_03632_),
    .B2(addr_i_2_),
    .Y(_08695_)
  );
  sg13g2_a22oi_1 _18360_ (
    .A1(addr_i_2_),
    .A2(_08694_),
    .B1(_08695_),
    .B2(_01674_),
    .Y(_08697_)
  );
  sg13g2_a21oi_1 _18361_ (
    .A1(_01441_),
    .A2(_01343_),
    .B1(addr_i_4_),
    .Y(_08698_)
  );
  sg13g2_or2_1 _18362_ (
    .A(_08697_),
    .B(_08698_),
    .X(_08699_)
  );
  sg13g2_o21ai_1 _18363_ (
    .A1(_08693_),
    .A2(_08699_),
    .B1(addr_i_8_),
    .Y(_08700_)
  );
  sg13g2_o21ai_1 _18364_ (
    .A1(_00607_),
    .A2(_01902_),
    .B1(addr_i_6_),
    .Y(_08701_)
  );
  sg13g2_a21oi_1 _18365_ (
    .A1(_02536_),
    .A2(_07557_),
    .B1(_04068_),
    .Y(_08702_)
  );
  sg13g2_a21o_1 _18366_ (
    .A1(_00831_),
    .A2(_00502_),
    .B1(addr_i_6_),
    .X(_08703_)
  );
  sg13g2_nor2_1 _18367_ (
    .A(addr_i_7_),
    .B(_03565_),
    .Y(_08704_)
  );
  sg13g2_a221oi_1 _18368_ (
    .A1(_08701_),
    .A2(_08702_),
    .B1(_08703_),
    .B2(_08704_),
    .C1(addr_i_8_),
    .Y(_08705_)
  );
  sg13g2_inv_1 _18369_ (
    .A(_08705_),
    .Y(_08706_)
  );
  sg13g2_a21oi_1 _18370_ (
    .A1(_08700_),
    .A2(_08706_),
    .B1(addr_i_9_),
    .Y(_08709_)
  );
  sg13g2_a22oi_1 _18371_ (
    .A1(addr_i_9_),
    .A2(_08689_),
    .B1(_08709_),
    .B2(addr_i_10_),
    .Y(_08710_)
  );
  sg13g2_nor2_1 _18372_ (
    .A(_00476_),
    .B(_00666_),
    .Y(_08711_)
  );
  sg13g2_a21oi_1 _18373_ (
    .A1(_03964_),
    .A2(_02694_),
    .B1(addr_i_3_),
    .Y(_08712_)
  );
  sg13g2_o21ai_1 _18374_ (
    .A1(_08711_),
    .A2(_08712_),
    .B1(addr_i_4_),
    .Y(_08713_)
  );
  sg13g2_a21oi_1 _18375_ (
    .A1(_06419_),
    .A2(_04538_),
    .B1(_02126_),
    .Y(_08714_)
  );
  sg13g2_o21ai_1 _18376_ (
    .A1(addr_i_4_),
    .A2(_08714_),
    .B1(_07790_),
    .Y(_08715_)
  );
  sg13g2_a21oi_1 _18377_ (
    .A1(_00343_),
    .A2(_00021_),
    .B1(_09061_),
    .Y(_08716_)
  );
  sg13g2_o21ai_1 _18378_ (
    .A1(addr_i_5_),
    .A2(_08716_),
    .B1(_01008_),
    .Y(_08717_)
  );
  sg13g2_o21ai_1 _18379_ (
    .A1(_03964_),
    .A2(_00697_),
    .B1(_03617_),
    .Y(_08718_)
  );
  sg13g2_a221oi_1 _18380_ (
    .A1(addr_i_2_),
    .A2(_08715_),
    .B1(_08717_),
    .B2(addr_i_3_),
    .C1(_08718_),
    .Y(_08720_)
  );
  sg13g2_a21oi_1 _18381_ (
    .A1(addr_i_7_),
    .A2(_00284_),
    .B1(_02479_),
    .Y(_08721_)
  );
  sg13g2_a22oi_1 _18382_ (
    .A1(_07248_),
    .A2(_02517_),
    .B1(_08721_),
    .B2(_00096_),
    .Y(_08722_)
  );
  sg13g2_a21oi_1 _18383_ (
    .A1(_04830_),
    .A2(_08722_),
    .B1(addr_i_3_),
    .Y(_08723_)
  );
  sg13g2_o21ai_1 _18384_ (
    .A1(_01114_),
    .A2(_02091_),
    .B1(_01301_),
    .Y(_08724_)
  );
  sg13g2_nand2_1 _18385_ (
    .A(addr_i_3_),
    .B(_04741_),
    .Y(_08725_)
  );
  sg13g2_nand2b_1 _18386_ (
    .A_N(_08725_),
    .B(_01950_),
    .Y(_08726_)
  );
  sg13g2_a21oi_1 _18387_ (
    .A1(_00146_),
    .A2(_08724_),
    .B1(_08726_),
    .Y(_08727_)
  );
  sg13g2_nor4_1 _18388_ (
    .A(_00782_),
    .B(_02542_),
    .C(_08723_),
    .D(_08727_),
    .Y(_08728_)
  );
  sg13g2_a21oi_1 _18389_ (
    .A1(_08713_),
    .A2(_08720_),
    .B1(_08728_),
    .Y(_08729_)
  );
  sg13g2_o21ai_1 _18390_ (
    .A1(_01070_),
    .A2(_05960_),
    .B1(_01290_),
    .Y(_08731_)
  );
  sg13g2_nand2_1 _18391_ (
    .A(_00380_),
    .B(_01273_),
    .Y(_08732_)
  );
  sg13g2_a22oi_1 _18392_ (
    .A1(addr_i_3_),
    .A2(_08732_),
    .B1(_02014_),
    .B2(_09359_),
    .Y(_08733_)
  );
  sg13g2_nor2_1 _18393_ (
    .A(addr_i_7_),
    .B(_08733_),
    .Y(_08734_)
  );
  sg13g2_a221oi_1 _18394_ (
    .A1(_04539_),
    .A2(_01065_),
    .B1(_07641_),
    .B2(_05402_),
    .C1(_01232_),
    .Y(_08735_)
  );
  sg13g2_a21oi_1 _18395_ (
    .A1(addr_i_7_),
    .A2(_00380_),
    .B1(_00120_),
    .Y(_08736_)
  );
  sg13g2_o21ai_1 _18396_ (
    .A1(_02238_),
    .A2(_08736_),
    .B1(_02777_),
    .Y(_08737_)
  );
  sg13g2_a21oi_1 _18397_ (
    .A1(_08735_),
    .A2(_08737_),
    .B1(addr_i_3_),
    .Y(_08738_)
  );
  sg13g2_a22oi_1 _18398_ (
    .A1(addr_i_3_),
    .A2(_08731_),
    .B1(_08734_),
    .B2(_08738_),
    .Y(_08739_)
  );
  sg13g2_nor2_1 _18399_ (
    .A(addr_i_8_),
    .B(_08739_),
    .Y(_08740_)
  );
  sg13g2_a21oi_1 _18400_ (
    .A1(_00147_),
    .A2(_01813_),
    .B1(addr_i_2_),
    .Y(_08742_)
  );
  sg13g2_o21ai_1 _18401_ (
    .A1(_01660_),
    .A2(_08742_),
    .B1(addr_i_7_),
    .Y(_08743_)
  );
  sg13g2_nand3_1 _18402_ (
    .A(_02683_),
    .B(_02047_),
    .C(_08743_),
    .Y(_08744_)
  );
  sg13g2_nor2_1 _18403_ (
    .A(addr_i_4_),
    .B(_01054_),
    .Y(_08745_)
  );
  sg13g2_o21ai_1 _18404_ (
    .A1(_03250_),
    .A2(_08745_),
    .B1(_01480_),
    .Y(_08746_)
  );
  sg13g2_a21o_1 _18405_ (
    .A1(_00994_),
    .A2(_00975_),
    .B1(_01514_),
    .X(_08747_)
  );
  sg13g2_nand3_1 _18406_ (
    .A(_05427_),
    .B(_08746_),
    .C(_08747_),
    .Y(_08748_)
  );
  sg13g2_a22oi_1 _18407_ (
    .A1(addr_i_3_),
    .A2(_08744_),
    .B1(_08748_),
    .B2(_01151_),
    .Y(_08749_)
  );
  sg13g2_nor3_1 _18408_ (
    .A(_00243_),
    .B(_08740_),
    .C(_08749_),
    .Y(_08750_)
  );
  sg13g2_a22oi_1 _18409_ (
    .A1(_00397_),
    .A2(_08729_),
    .B1(_08750_),
    .B2(_01774_),
    .Y(_08751_)
  );
  sg13g2_o21ai_1 _18410_ (
    .A1(_08710_),
    .A2(_08751_),
    .B1(_03051_),
    .Y(_08753_)
  );
  sg13g2_a21o_1 _18411_ (
    .A1(addr_i_3_),
    .A2(_02948_),
    .B1(_01107_),
    .X(_08754_)
  );
  sg13g2_o21ai_1 _18412_ (
    .A1(addr_i_4_),
    .A2(_03245_),
    .B1(_01067_),
    .Y(_08755_)
  );
  sg13g2_a21oi_1 _18413_ (
    .A1(_01029_),
    .A2(_08755_),
    .B1(addr_i_5_),
    .Y(_08756_)
  );
  sg13g2_a22oi_1 _18414_ (
    .A1(addr_i_6_),
    .A2(_08754_),
    .B1(_08756_),
    .B2(addr_i_7_),
    .Y(_08757_)
  );
  sg13g2_nor2_1 _18415_ (
    .A(_00645_),
    .B(_08757_),
    .Y(_08758_)
  );
  sg13g2_o21ai_1 _18416_ (
    .A1(_01007_),
    .A2(_01486_),
    .B1(_01343_),
    .Y(_08759_)
  );
  sg13g2_nand2_1 _18417_ (
    .A(addr_i_3_),
    .B(_00477_),
    .Y(_08760_)
  );
  sg13g2_a22oi_1 _18418_ (
    .A1(_02012_),
    .A2(_08760_),
    .B1(_00083_),
    .B2(addr_i_7_),
    .Y(_08761_)
  );
  sg13g2_a21oi_1 _18419_ (
    .A1(_02803_),
    .A2(_08759_),
    .B1(_08761_),
    .Y(_08762_)
  );
  sg13g2_nand2_1 _18420_ (
    .A(_00573_),
    .B(_03324_),
    .Y(_08764_)
  );
  sg13g2_a21oi_1 _18421_ (
    .A1(_02930_),
    .A2(_00453_),
    .B1(addr_i_3_),
    .Y(_08765_)
  );
  sg13g2_a21oi_1 _18422_ (
    .A1(_02470_),
    .A2(_00668_),
    .B1(addr_i_5_),
    .Y(_08766_)
  );
  sg13g2_a22oi_1 _18423_ (
    .A1(addr_i_7_),
    .A2(_08764_),
    .B1(_08765_),
    .B2(_08766_),
    .Y(_08767_)
  );
  sg13g2_a21oi_1 _18424_ (
    .A1(_08762_),
    .A2(_08767_),
    .B1(addr_i_8_),
    .Y(_08768_)
  );
  sg13g2_a22oi_1 _18425_ (
    .A1(addr_i_8_),
    .A2(_08758_),
    .B1(_08768_),
    .B2(addr_i_9_),
    .Y(_08769_)
  );
  sg13g2_nor2b_1 _18426_ (
    .A(_08769_),
    .B_N(_05074_),
    .Y(_08770_)
  );
  sg13g2_a22oi_1 _18427_ (
    .A1(_03084_),
    .A2(_03829_),
    .B1(_05099_),
    .B2(_08770_),
    .Y(_08771_)
  );
  sg13g2_nor2_1 _18428_ (
    .A(_00812_),
    .B(_08771_),
    .Y(_08772_)
  );
  sg13g2_nand2_1 _18429_ (
    .A(_05025_),
    .B(_00665_),
    .Y(_08773_)
  );
  sg13g2_o21ai_1 _18430_ (
    .A1(_00543_),
    .A2(_02761_),
    .B1(_08773_),
    .Y(_08775_)
  );
  sg13g2_a221oi_1 _18431_ (
    .A1(_08598_),
    .A2(_00301_),
    .B1(_08775_),
    .B2(addr_i_2_),
    .C1(addr_i_8_),
    .Y(_08776_)
  );
  sg13g2_o21ai_1 _18432_ (
    .A1(_00581_),
    .A2(_00194_),
    .B1(_04395_),
    .Y(_08777_)
  );
  sg13g2_nand2_1 _18433_ (
    .A(_06607_),
    .B(_08777_),
    .Y(_08778_)
  );
  sg13g2_a21o_1 _18434_ (
    .A1(_04741_),
    .A2(_08778_),
    .B1(addr_i_3_),
    .X(_08779_)
  );
  sg13g2_a21oi_1 _18435_ (
    .A1(_01120_),
    .A2(_02405_),
    .B1(_02153_),
    .Y(_08780_)
  );
  sg13g2_nor2_1 _18436_ (
    .A(addr_i_2_),
    .B(_08780_),
    .Y(_08781_)
  );
  sg13g2_o21ai_1 _18437_ (
    .A1(_02479_),
    .A2(_01658_),
    .B1(_06292_),
    .Y(_08782_)
  );
  sg13g2_o21ai_1 _18438_ (
    .A1(_08781_),
    .A2(_08782_),
    .B1(addr_i_3_),
    .Y(_08783_)
  );
  sg13g2_nand3_1 _18439_ (
    .A(_08776_),
    .B(_08779_),
    .C(_08783_),
    .Y(_08784_)
  );
  sg13g2_o21ai_1 _18440_ (
    .A1(_04108_),
    .A2(_01507_),
    .B1(_02349_),
    .Y(_08786_)
  );
  sg13g2_a21oi_1 _18441_ (
    .A1(_08707_),
    .A2(_02822_),
    .B1(_08000_),
    .Y(_08787_)
  );
  sg13g2_a22oi_1 _18442_ (
    .A1(_05867_),
    .A2(_08786_),
    .B1(_08787_),
    .B2(_00227_),
    .Y(_08788_)
  );
  sg13g2_a22oi_1 _18443_ (
    .A1(addr_i_4_),
    .A2(_00736_),
    .B1(_00597_),
    .B2(_00059_),
    .Y(_08789_)
  );
  sg13g2_a22oi_1 _18444_ (
    .A1(_09491_),
    .A2(_02725_),
    .B1(_08789_),
    .B2(addr_i_7_),
    .Y(_08790_)
  );
  sg13g2_nor2_1 _18445_ (
    .A(_07282_),
    .B(_08790_),
    .Y(_08791_)
  );
  sg13g2_o21ai_1 _18446_ (
    .A1(_04052_),
    .A2(_08788_),
    .B1(_08791_),
    .Y(_08792_)
  );
  sg13g2_nand3_1 _18447_ (
    .A(_01351_),
    .B(_08784_),
    .C(_08792_),
    .Y(_08793_)
  );
  sg13g2_o21ai_1 _18448_ (
    .A1(_07359_),
    .A2(_00635_),
    .B1(addr_i_2_),
    .Y(_08794_)
  );
  sg13g2_mux2_1 _18449_ (
    .A0(_07222_),
    .A1(_07943_),
    .S(_08156_),
    .X(_08795_)
  );
  sg13g2_a21oi_1 _18450_ (
    .A1(_08794_),
    .A2(_08795_),
    .B1(addr_i_5_),
    .Y(_08797_)
  );
  sg13g2_a21oi_1 _18451_ (
    .A1(_00117_),
    .A2(_08929_),
    .B1(addr_i_6_),
    .Y(_08798_)
  );
  sg13g2_a21oi_1 _18452_ (
    .A1(_01579_),
    .A2(_04747_),
    .B1(_08798_),
    .Y(_08799_)
  );
  sg13g2_a21oi_1 _18453_ (
    .A1(_04151_),
    .A2(_01319_),
    .B1(addr_i_8_),
    .Y(_08800_)
  );
  sg13g2_o21ai_1 _18454_ (
    .A1(addr_i_2_),
    .A2(_08799_),
    .B1(_08800_),
    .Y(_08801_)
  );
  sg13g2_o21ai_1 _18455_ (
    .A1(_08797_),
    .A2(_08801_),
    .B1(addr_i_9_),
    .Y(_08802_)
  );
  sg13g2_o21ai_1 _18456_ (
    .A1(_00269_),
    .A2(_01375_),
    .B1(_09127_),
    .Y(_08803_)
  );
  sg13g2_a21oi_1 _18457_ (
    .A1(_09497_),
    .A2(_02200_),
    .B1(_00010_),
    .Y(_08804_)
  );
  sg13g2_a21oi_1 _18458_ (
    .A1(_08803_),
    .A2(_08804_),
    .B1(addr_i_3_),
    .Y(_08805_)
  );
  sg13g2_a21oi_1 _18459_ (
    .A1(_02349_),
    .A2(_09371_),
    .B1(addr_i_4_),
    .Y(_08806_)
  );
  sg13g2_a22oi_1 _18460_ (
    .A1(_09127_),
    .A2(_08144_),
    .B1(_01112_),
    .B2(_08806_),
    .Y(_08808_)
  );
  sg13g2_nor3_1 _18461_ (
    .A(_00535_),
    .B(addr_i_4_),
    .C(_01054_),
    .Y(_08809_)
  );
  sg13g2_a21oi_1 _18462_ (
    .A1(_00016_),
    .A2(_00973_),
    .B1(_00956_),
    .Y(_08810_)
  );
  sg13g2_o21ai_1 _18463_ (
    .A1(_08809_),
    .A2(_08810_),
    .B1(_00200_),
    .Y(_08811_)
  );
  sg13g2_o21ai_1 _18464_ (
    .A1(_00799_),
    .A2(_08808_),
    .B1(_08811_),
    .Y(_08812_)
  );
  sg13g2_o21ai_1 _18465_ (
    .A1(_08805_),
    .A2(_08812_),
    .B1(addr_i_8_),
    .Y(_08813_)
  );
  sg13g2_nand2b_1 _18466_ (
    .A_N(_08802_),
    .B(_08813_),
    .Y(_08814_)
  );
  sg13g2_a21oi_1 _18467_ (
    .A1(_08793_),
    .A2(_08814_),
    .B1(_03841_),
    .Y(_08815_)
  );
  sg13g2_o21ai_1 _18468_ (
    .A1(_05014_),
    .A2(_05524_),
    .B1(addr_i_3_),
    .Y(_08816_)
  );
  sg13g2_nand3_1 _18469_ (
    .A(_04087_),
    .B(_02136_),
    .C(_08816_),
    .Y(_08817_)
  );
  sg13g2_a22oi_1 _18470_ (
    .A1(addr_i_5_),
    .A2(_08817_),
    .B1(_05005_),
    .B2(_07951_),
    .Y(_08820_)
  );
  sg13g2_nand2_1 _18471_ (
    .A(_00831_),
    .B(_00649_),
    .Y(_08821_)
  );
  sg13g2_o21ai_1 _18472_ (
    .A1(_03648_),
    .A2(_01791_),
    .B1(addr_i_8_),
    .Y(_08822_)
  );
  sg13g2_nor4_1 _18473_ (
    .A(_02569_),
    .B(_06795_),
    .C(_03033_),
    .D(_03846_),
    .Y(_08823_)
  );
  sg13g2_a22oi_1 _18474_ (
    .A1(_01320_),
    .A2(_08821_),
    .B1(_08822_),
    .B2(_08823_),
    .Y(_08824_)
  );
  sg13g2_o21ai_1 _18475_ (
    .A1(_02257_),
    .A2(_08820_),
    .B1(_08824_),
    .Y(_08825_)
  );
  sg13g2_mux2_1 _18476_ (
    .A0(_00086_),
    .A1(_00210_),
    .S(addr_i_5_),
    .X(_08826_)
  );
  sg13g2_a21oi_1 _18477_ (
    .A1(addr_i_7_),
    .A2(_00024_),
    .B1(addr_i_3_),
    .Y(_08827_)
  );
  sg13g2_a21oi_1 _18478_ (
    .A1(addr_i_4_),
    .A2(_08826_),
    .B1(_08827_),
    .Y(_08828_)
  );
  sg13g2_a21oi_1 _18479_ (
    .A1(_01603_),
    .A2(_00680_),
    .B1(_03864_),
    .Y(_08829_)
  );
  sg13g2_o21ai_1 _18480_ (
    .A1(_01127_),
    .A2(_08829_),
    .B1(addr_i_4_),
    .Y(_08831_)
  );
  sg13g2_o21ai_1 _18481_ (
    .A1(_04251_),
    .A2(_08828_),
    .B1(_08831_),
    .Y(_08832_)
  );
  sg13g2_nand3_1 _18482_ (
    .A(_00091_),
    .B(_00294_),
    .C(_01208_),
    .Y(_08833_)
  );
  sg13g2_nor3_1 _18483_ (
    .A(_02086_),
    .B(addr_i_5_),
    .C(_05236_),
    .Y(_08834_)
  );
  sg13g2_o21ai_1 _18484_ (
    .A1(_03793_),
    .A2(_08834_),
    .B1(_00145_),
    .Y(_08835_)
  );
  sg13g2_a21oi_1 _18485_ (
    .A1(_08833_),
    .A2(_08835_),
    .B1(addr_i_4_),
    .Y(_08836_)
  );
  sg13g2_o21ai_1 _18486_ (
    .A1(_08832_),
    .A2(_08836_),
    .B1(_01043_),
    .Y(_08837_)
  );
  sg13g2_nand3_1 _18487_ (
    .A(addr_i_9_),
    .B(_08825_),
    .C(_08837_),
    .Y(_08838_)
  );
  sg13g2_nand2_1 _18488_ (
    .A(_00020_),
    .B(_03424_),
    .Y(_08839_)
  );
  sg13g2_o21ai_1 _18489_ (
    .A1(_01252_),
    .A2(_01495_),
    .B1(_01912_),
    .Y(_08840_)
  );
  sg13g2_nor2_1 _18490_ (
    .A(addr_i_6_),
    .B(_02448_),
    .Y(_08842_)
  );
  sg13g2_a22oi_1 _18491_ (
    .A1(_06806_),
    .A2(_08839_),
    .B1(_08840_),
    .B2(_08842_),
    .Y(_08843_)
  );
  sg13g2_a21o_1 _18492_ (
    .A1(addr_i_4_),
    .A2(_01486_),
    .B1(_00247_),
    .X(_08844_)
  );
  sg13g2_a21o_1 _18493_ (
    .A1(_02031_),
    .A2(_00926_),
    .B1(_03864_),
    .X(_08845_)
  );
  sg13g2_o21ai_1 _18494_ (
    .A1(_00052_),
    .A2(_02536_),
    .B1(_08845_),
    .Y(_08846_)
  );
  sg13g2_a221oi_1 _18495_ (
    .A1(_03348_),
    .A2(_08844_),
    .B1(_08846_),
    .B2(_08708_),
    .C1(_07282_),
    .Y(_08847_)
  );
  sg13g2_o21ai_1 _18496_ (
    .A1(addr_i_3_),
    .A2(_08843_),
    .B1(_08847_),
    .Y(_08848_)
  );
  sg13g2_a21oi_1 _18497_ (
    .A1(_01603_),
    .A2(_01729_),
    .B1(_09491_),
    .Y(_08849_)
  );
  sg13g2_o21ai_1 _18498_ (
    .A1(_00945_),
    .A2(_08849_),
    .B1(addr_i_4_),
    .Y(_08850_)
  );
  sg13g2_a221oi_1 _18499_ (
    .A1(_05689_),
    .A2(_00583_),
    .B1(_05746_),
    .B2(_01033_),
    .C1(_05070_),
    .Y(_08851_)
  );
  sg13g2_a22oi_1 _18500_ (
    .A1(_00483_),
    .A2(_00184_),
    .B1(_03139_),
    .B2(addr_i_7_),
    .Y(_08853_)
  );
  sg13g2_nor2_1 _18501_ (
    .A(_08851_),
    .B(_08853_),
    .Y(_08854_)
  );
  sg13g2_nor2_1 _18502_ (
    .A(addr_i_8_),
    .B(_08854_),
    .Y(_08855_)
  );
  sg13g2_a21oi_1 _18503_ (
    .A1(_08850_),
    .A2(_08855_),
    .B1(addr_i_9_),
    .Y(_08856_)
  );
  sg13g2_a21oi_1 _18504_ (
    .A1(_08848_),
    .A2(_08856_),
    .B1(addr_i_10_),
    .Y(_08857_)
  );
  sg13g2_a21oi_1 _18505_ (
    .A1(_08838_),
    .A2(_08857_),
    .B1(addr_i_11_),
    .Y(_08858_)
  );
  sg13g2_nand2b_1 _18506_ (
    .A_N(_08815_),
    .B(_08858_),
    .Y(_08859_)
  );
  sg13g2_a22oi_1 _18507_ (
    .A1(_00044_),
    .A2(_05225_),
    .B1(_05014_),
    .B2(_00064_),
    .Y(_08860_)
  );
  sg13g2_or2_1 _18508_ (
    .A(_07215_),
    .B(_08860_),
    .X(_08861_)
  );
  sg13g2_a22oi_1 _18509_ (
    .A1(addr_i_5_),
    .A2(_00254_),
    .B1(_07998_),
    .B2(_06607_),
    .Y(_08862_)
  );
  sg13g2_a21oi_1 _18510_ (
    .A1(_00200_),
    .A2(_08861_),
    .B1(_08862_),
    .Y(_08864_)
  );
  sg13g2_o21ai_1 _18511_ (
    .A1(_00914_),
    .A2(_00304_),
    .B1(_02440_),
    .Y(_08865_)
  );
  sg13g2_o21ai_1 _18512_ (
    .A1(_00679_),
    .A2(_00304_),
    .B1(_00863_),
    .Y(_08866_)
  );
  sg13g2_a22oi_1 _18513_ (
    .A1(addr_i_7_),
    .A2(_08865_),
    .B1(_08866_),
    .B2(addr_i_3_),
    .Y(_08867_)
  );
  sg13g2_a22oi_1 _18514_ (
    .A1(addr_i_3_),
    .A2(_08864_),
    .B1(_08867_),
    .B2(addr_i_8_),
    .Y(_08868_)
  );
  sg13g2_a22oi_1 _18515_ (
    .A1(_01652_),
    .A2(_00686_),
    .B1(_03416_),
    .B2(addr_i_4_),
    .Y(_08869_)
  );
  sg13g2_nand3_1 _18516_ (
    .A(addr_i_4_),
    .B(_00050_),
    .C(_07624_),
    .Y(_08870_)
  );
  sg13g2_nor2b_1 _18517_ (
    .A(_08869_),
    .B_N(_08870_),
    .Y(_08871_)
  );
  sg13g2_o21ai_1 _18518_ (
    .A1(_01436_),
    .A2(_05634_),
    .B1(addr_i_3_),
    .Y(_08872_)
  );
  sg13g2_nor3_1 _18519_ (
    .A(_06496_),
    .B(_00165_),
    .C(_00521_),
    .Y(_08873_)
  );
  sg13g2_a221oi_1 _18520_ (
    .A1(_04284_),
    .A2(_01652_),
    .B1(_01436_),
    .B2(_08376_),
    .C1(_08873_),
    .Y(_08875_)
  );
  sg13g2_a21oi_1 _18521_ (
    .A1(_08872_),
    .A2(_08875_),
    .B1(addr_i_2_),
    .Y(_08876_)
  );
  sg13g2_o21ai_1 _18522_ (
    .A1(_08871_),
    .A2(_08876_),
    .B1(addr_i_8_),
    .Y(_08877_)
  );
  sg13g2_nand2b_1 _18523_ (
    .A_N(_08868_),
    .B(_08877_),
    .Y(_08878_)
  );
  sg13g2_a22oi_1 _18524_ (
    .A1(addr_i_4_),
    .A2(_04854_),
    .B1(_01604_),
    .B2(addr_i_8_),
    .Y(_08879_)
  );
  sg13g2_o21ai_1 _18525_ (
    .A1(_00294_),
    .A2(_01867_),
    .B1(addr_i_4_),
    .Y(_08880_)
  );
  sg13g2_o21ai_1 _18526_ (
    .A1(_03776_),
    .A2(_00384_),
    .B1(_00065_),
    .Y(_08881_)
  );
  sg13g2_nand3_1 _18527_ (
    .A(_03258_),
    .B(_08880_),
    .C(_08881_),
    .Y(_08882_)
  );
  sg13g2_nand3_1 _18528_ (
    .A(_00927_),
    .B(_03540_),
    .C(_07359_),
    .Y(_08883_)
  );
  sg13g2_o21ai_1 _18529_ (
    .A1(_00977_),
    .A2(_05634_),
    .B1(addr_i_4_),
    .Y(_08884_)
  );
  sg13g2_nand4_1 _18530_ (
    .A(addr_i_3_),
    .B(_04295_),
    .C(_08883_),
    .D(_08884_),
    .Y(_08886_)
  );
  sg13g2_o21ai_1 _18531_ (
    .A1(addr_i_3_),
    .A2(_08882_),
    .B1(_08886_),
    .Y(_08887_)
  );
  sg13g2_o21ai_1 _18532_ (
    .A1(_09513_),
    .A2(_02732_),
    .B1(_01921_),
    .Y(_08888_)
  );
  sg13g2_nor2_1 _18533_ (
    .A(addr_i_3_),
    .B(_00376_),
    .Y(_08889_)
  );
  sg13g2_nor2_1 _18534_ (
    .A(_04981_),
    .B(_06752_),
    .Y(_08890_)
  );
  sg13g2_a22oi_1 _18535_ (
    .A1(_08232_),
    .A2(_08889_),
    .B1(_08890_),
    .B2(_00949_),
    .Y(_08891_)
  );
  sg13g2_nor3_1 _18536_ (
    .A(_00297_),
    .B(_08144_),
    .C(_02107_),
    .Y(_08892_)
  );
  sg13g2_a21oi_1 _18537_ (
    .A1(_00566_),
    .A2(_03267_),
    .B1(_06684_),
    .Y(_08893_)
  );
  sg13g2_o21ai_1 _18538_ (
    .A1(addr_i_6_),
    .A2(_08892_),
    .B1(_08893_),
    .Y(_08894_)
  );
  sg13g2_a22oi_1 _18539_ (
    .A1(_05822_),
    .A2(_08888_),
    .B1(_08891_),
    .B2(_08894_),
    .Y(_08895_)
  );
  sg13g2_a22oi_1 _18540_ (
    .A1(_08879_),
    .A2(_08887_),
    .B1(_08895_),
    .B2(addr_i_9_),
    .Y(_08897_)
  );
  sg13g2_a22oi_1 _18541_ (
    .A1(addr_i_9_),
    .A2(_08878_),
    .B1(_08897_),
    .B2(_01773_),
    .Y(_08898_)
  );
  sg13g2_o21ai_1 _18542_ (
    .A1(_00199_),
    .A2(_07871_),
    .B1(_01029_),
    .Y(_08899_)
  );
  sg13g2_a21oi_1 _18543_ (
    .A1(_00435_),
    .A2(_02031_),
    .B1(addr_i_5_),
    .Y(_08900_)
  );
  sg13g2_a22oi_1 _18544_ (
    .A1(addr_i_7_),
    .A2(_08899_),
    .B1(_08900_),
    .B2(_03137_),
    .Y(_08901_)
  );
  sg13g2_nand2b_1 _18545_ (
    .A_N(_08901_),
    .B(addr_i_3_),
    .Y(_08902_)
  );
  sg13g2_o21ai_1 _18546_ (
    .A1(addr_i_2_),
    .A2(_07027_),
    .B1(_01658_),
    .Y(_08903_)
  );
  sg13g2_a21oi_1 _18547_ (
    .A1(_04804_),
    .A2(_03875_),
    .B1(addr_i_5_),
    .Y(_08904_)
  );
  sg13g2_a21o_1 _18548_ (
    .A1(_08785_),
    .A2(_08903_),
    .B1(_08904_),
    .X(_08905_)
  );
  sg13g2_a21oi_1 _18549_ (
    .A1(_00434_),
    .A2(_00037_),
    .B1(_00104_),
    .Y(_08906_)
  );
  sg13g2_o21ai_1 _18550_ (
    .A1(_00692_),
    .A2(_02089_),
    .B1(addr_i_8_),
    .Y(_08908_)
  );
  sg13g2_a22oi_1 _18551_ (
    .A1(addr_i_4_),
    .A2(_08905_),
    .B1(_08906_),
    .B2(_08908_),
    .Y(_08909_)
  );
  sg13g2_o21ai_1 _18552_ (
    .A1(_02634_),
    .A2(_00448_),
    .B1(_01175_),
    .Y(_08910_)
  );
  sg13g2_a21oi_1 _18553_ (
    .A1(_00550_),
    .A2(_08852_),
    .B1(_00780_),
    .Y(_08911_)
  );
  sg13g2_nand2_1 _18554_ (
    .A(_02434_),
    .B(_08911_),
    .Y(_08912_)
  );
  sg13g2_a221oi_1 _18555_ (
    .A1(_01355_),
    .A2(_02166_),
    .B1(_08910_),
    .B2(_00726_),
    .C1(_08912_),
    .Y(_08913_)
  );
  sg13g2_nor2_1 _18556_ (
    .A(_05402_),
    .B(_00334_),
    .Y(_08914_)
  );
  sg13g2_nand2_1 _18557_ (
    .A(_04981_),
    .B(_06790_),
    .Y(_08915_)
  );
  sg13g2_a21oi_1 _18558_ (
    .A1(addr_i_3_),
    .A2(_00665_),
    .B1(addr_i_4_),
    .Y(_08916_)
  );
  sg13g2_a221oi_1 _18559_ (
    .A1(_07542_),
    .A2(_08914_),
    .B1(_08915_),
    .B2(_08916_),
    .C1(_07603_),
    .Y(_08917_)
  );
  sg13g2_a22oi_1 _18560_ (
    .A1(_08902_),
    .A2(_08909_),
    .B1(_08913_),
    .B2(_08917_),
    .Y(_08919_)
  );
  sg13g2_nand2b_1 _18561_ (
    .A_N(_08919_),
    .B(addr_i_9_),
    .Y(_08920_)
  );
  sg13g2_o21ai_1 _18562_ (
    .A1(_02055_),
    .A2(_06271_),
    .B1(addr_i_3_),
    .Y(_08921_)
  );
  sg13g2_nand2_1 _18563_ (
    .A(_00651_),
    .B(_05964_),
    .Y(_08922_)
  );
  sg13g2_a21oi_1 _18564_ (
    .A1(_02810_),
    .A2(_00870_),
    .B1(_02796_),
    .Y(_08923_)
  );
  sg13g2_a22oi_1 _18565_ (
    .A1(_02257_),
    .A2(_08922_),
    .B1(_08923_),
    .B2(_03494_),
    .Y(_08924_)
  );
  sg13g2_nand2_1 _18566_ (
    .A(_08921_),
    .B(_08924_),
    .Y(_08925_)
  );
  sg13g2_o21ai_1 _18567_ (
    .A1(_08653_),
    .A2(_01571_),
    .B1(_00083_),
    .Y(_08926_)
  );
  sg13g2_nand3_1 _18568_ (
    .A(addr_i_3_),
    .B(_00148_),
    .C(_05318_),
    .Y(_08927_)
  );
  sg13g2_o21ai_1 _18569_ (
    .A1(addr_i_3_),
    .A2(_08546_),
    .B1(_08927_),
    .Y(_08928_)
  );
  sg13g2_a21oi_1 _18570_ (
    .A1(_08926_),
    .A2(_08928_),
    .B1(_02963_),
    .Y(_08931_)
  );
  sg13g2_a21oi_1 _18571_ (
    .A1(addr_i_3_),
    .A2(_00520_),
    .B1(_02297_),
    .Y(_08932_)
  );
  sg13g2_nand2_1 _18572_ (
    .A(addr_i_3_),
    .B(_01813_),
    .Y(_08933_)
  );
  sg13g2_a21oi_1 _18573_ (
    .A1(_05613_),
    .A2(_08933_),
    .B1(_02344_),
    .Y(_08934_)
  );
  sg13g2_nor4_1 _18574_ (
    .A(_00206_),
    .B(_03203_),
    .C(_08932_),
    .D(_08934_),
    .Y(_08935_)
  );
  sg13g2_o21ai_1 _18575_ (
    .A1(_00726_),
    .A2(_06088_),
    .B1(_08431_),
    .Y(_08936_)
  );
  sg13g2_nand2_1 _18576_ (
    .A(_09491_),
    .B(_04077_),
    .Y(_08937_)
  );
  sg13g2_a21oi_1 _18577_ (
    .A1(_04866_),
    .A2(_08937_),
    .B1(_00067_),
    .Y(_08938_)
  );
  sg13g2_a22oi_1 _18578_ (
    .A1(_00818_),
    .A2(_08936_),
    .B1(_08938_),
    .B2(_02535_),
    .Y(_08939_)
  );
  sg13g2_nor4_1 _18579_ (
    .A(addr_i_10_),
    .B(_08931_),
    .C(_08935_),
    .D(_08939_),
    .Y(_08940_)
  );
  sg13g2_nand3_1 _18580_ (
    .A(_08920_),
    .B(_08925_),
    .C(_08940_),
    .Y(_08942_)
  );
  sg13g2_nand3b_1 _18581_ (
    .A_N(_08898_),
    .B(_08942_),
    .C(addr_i_11_),
    .Y(_08943_)
  );
  sg13g2_a21oi_1 _18582_ (
    .A1(_08859_),
    .A2(_08943_),
    .B1(addr_i_12_),
    .Y(_08944_)
  );
  sg13g2_a21o_1 _18583_ (
    .A1(_08753_),
    .A2(_08772_),
    .B1(_08944_),
    .X(data_o_7_)
  );
  sg13g2_o21ai_1 _18584_ (
    .A1(_00177_),
    .A2(_05361_),
    .B1(_02796_),
    .Y(_08945_)
  );
  sg13g2_a21oi_1 _18585_ (
    .A1(addr_i_2_),
    .A2(_00544_),
    .B1(_09494_),
    .Y(_08946_)
  );
  sg13g2_a21oi_1 _18586_ (
    .A1(_01108_),
    .A2(_08946_),
    .B1(_02759_),
    .Y(_08947_)
  );
  sg13g2_a21oi_1 _18587_ (
    .A1(_09513_),
    .A2(_00840_),
    .B1(_08653_),
    .Y(_08948_)
  );
  sg13g2_o21ai_1 _18588_ (
    .A1(_00548_),
    .A2(_08948_),
    .B1(addr_i_8_),
    .Y(_08949_)
  );
  sg13g2_a22oi_1 _18589_ (
    .A1(_08704_),
    .A2(_08945_),
    .B1(_08947_),
    .B2(_08949_),
    .Y(_08950_)
  );
  sg13g2_a22oi_1 _18590_ (
    .A1(_00072_),
    .A2(_08410_),
    .B1(_08575_),
    .B2(_01016_),
    .Y(_08952_)
  );
  sg13g2_nand2_1 _18591_ (
    .A(_00284_),
    .B(_01353_),
    .Y(_08953_)
  );
  sg13g2_a22oi_1 _18592_ (
    .A1(_01355_),
    .A2(_08953_),
    .B1(addr_i_8_),
    .B2(_00587_),
    .Y(_08954_)
  );
  sg13g2_o21ai_1 _18593_ (
    .A1(_03263_),
    .A2(_08952_),
    .B1(_08954_),
    .Y(_08955_)
  );
  sg13g2_a22oi_1 _18594_ (
    .A1(addr_i_3_),
    .A2(_02943_),
    .B1(_02500_),
    .B2(_00899_),
    .Y(_08956_)
  );
  sg13g2_a21oi_1 _18595_ (
    .A1(_00802_),
    .A2(_08955_),
    .B1(_08956_),
    .Y(_08957_)
  );
  sg13g2_nor2_1 _18596_ (
    .A(_08950_),
    .B(_08957_),
    .Y(_08958_)
  );
  sg13g2_nor4_1 _18597_ (
    .A(_01365_),
    .B(_01787_),
    .C(_02179_),
    .D(_02925_),
    .Y(_08959_)
  );
  sg13g2_o21ai_1 _18598_ (
    .A1(_08958_),
    .A2(_08959_),
    .B1(_01176_),
    .Y(_08960_)
  );
  sg13g2_o21ai_1 _18599_ (
    .A1(addr_i_3_),
    .A2(_05960_),
    .B1(_07177_),
    .Y(_08961_)
  );
  sg13g2_nor3_1 _18600_ (
    .A(_00338_),
    .B(_02055_),
    .C(_08961_),
    .Y(_08963_)
  );
  sg13g2_a22oi_1 _18601_ (
    .A1(_00838_),
    .A2(_03077_),
    .B1(_00794_),
    .B2(_01285_),
    .Y(_08964_)
  );
  sg13g2_a21oi_1 _18602_ (
    .A1(addr_i_3_),
    .A2(_00118_),
    .B1(_00261_),
    .Y(_08965_)
  );
  sg13g2_nand2_1 _18603_ (
    .A(_07816_),
    .B(_08965_),
    .Y(_08966_)
  );
  sg13g2_o21ai_1 _18604_ (
    .A1(_06088_),
    .A2(_00244_),
    .B1(_02191_),
    .Y(_08967_)
  );
  sg13g2_a21oi_1 _18605_ (
    .A1(_07790_),
    .A2(_00943_),
    .B1(_00080_),
    .Y(_08968_)
  );
  sg13g2_a22oi_1 _18606_ (
    .A1(_01169_),
    .A2(_08967_),
    .B1(_08968_),
    .B2(_02562_),
    .Y(_08969_)
  );
  sg13g2_o21ai_1 _18607_ (
    .A1(_00840_),
    .A2(_03864_),
    .B1(_07790_),
    .Y(_08970_)
  );
  sg13g2_a22oi_1 _18608_ (
    .A1(addr_i_4_),
    .A2(_08970_),
    .B1(_02010_),
    .B2(_00600_),
    .Y(_08971_)
  );
  sg13g2_a22oi_1 _18609_ (
    .A1(_08964_),
    .A2(_08966_),
    .B1(_08969_),
    .B2(_08971_),
    .Y(_08972_)
  );
  sg13g2_o21ai_1 _18610_ (
    .A1(_03062_),
    .A2(_08963_),
    .B1(_08972_),
    .Y(_08974_)
  );
  sg13g2_a21oi_1 _18611_ (
    .A1(_05203_),
    .A2(_08974_),
    .B1(addr_i_11_),
    .Y(_08975_)
  );
  sg13g2_nand2_1 _18612_ (
    .A(_08960_),
    .B(_08975_),
    .Y(_08976_)
  );
  sg13g2_a21oi_1 _18613_ (
    .A1(addr_i_6_),
    .A2(_00927_),
    .B1(_08000_),
    .Y(_08977_)
  );
  sg13g2_nand3_1 _18614_ (
    .A(addr_i_3_),
    .B(_00405_),
    .C(_01004_),
    .Y(_08978_)
  );
  sg13g2_o21ai_1 _18615_ (
    .A1(addr_i_3_),
    .A2(_08977_),
    .B1(_08978_),
    .Y(_08979_)
  );
  sg13g2_nand2b_1 _18616_ (
    .A_N(_00023_),
    .B(_08979_),
    .Y(_08980_)
  );
  sg13g2_o21ai_1 _18617_ (
    .A1(_00069_),
    .A2(_07558_),
    .B1(_00507_),
    .Y(_08981_)
  );
  sg13g2_a21oi_1 _18618_ (
    .A1(addr_i_6_),
    .A2(_01603_),
    .B1(addr_i_5_),
    .Y(_08982_)
  );
  sg13g2_a221oi_1 _18619_ (
    .A1(_02742_),
    .A2(_02134_),
    .B1(_05746_),
    .B2(_06740_),
    .C1(_08982_),
    .Y(_08983_)
  );
  sg13g2_nor2_1 _18620_ (
    .A(addr_i_4_),
    .B(_08983_),
    .Y(_08985_)
  );
  sg13g2_a22oi_1 _18621_ (
    .A1(addr_i_4_),
    .A2(_08980_),
    .B1(_08981_),
    .B2(_08985_),
    .Y(_08986_)
  );
  sg13g2_nor3_1 _18622_ (
    .A(_00227_),
    .B(_03186_),
    .C(_01187_),
    .Y(_08987_)
  );
  sg13g2_o21ai_1 _18623_ (
    .A1(_00507_),
    .A2(_08987_),
    .B1(addr_i_8_),
    .Y(_08988_)
  );
  sg13g2_o21ai_1 _18624_ (
    .A1(_00297_),
    .A2(_02322_),
    .B1(_00861_),
    .Y(_08989_)
  );
  sg13g2_o21ai_1 _18625_ (
    .A1(_04539_),
    .A2(_02015_),
    .B1(addr_i_7_),
    .Y(_08990_)
  );
  sg13g2_nand3_1 _18626_ (
    .A(_02987_),
    .B(_08989_),
    .C(_08990_),
    .Y(_08991_)
  );
  sg13g2_o21ai_1 _18627_ (
    .A1(_02514_),
    .A2(_00278_),
    .B1(addr_i_4_),
    .Y(_08992_)
  );
  sg13g2_nand3_1 _18628_ (
    .A(_01104_),
    .B(_08533_),
    .C(_08992_),
    .Y(_08993_)
  );
  sg13g2_nand3_1 _18629_ (
    .A(_00262_),
    .B(_00651_),
    .C(_00314_),
    .Y(_08994_)
  );
  sg13g2_nand2_1 _18630_ (
    .A(_06695_),
    .B(_08994_),
    .Y(_08996_)
  );
  sg13g2_a221oi_1 _18631_ (
    .A1(addr_i_6_),
    .A2(_08991_),
    .B1(_08993_),
    .B2(_01542_),
    .C1(_08996_),
    .Y(_08997_)
  );
  sg13g2_nor2_1 _18632_ (
    .A(_00396_),
    .B(_08997_),
    .Y(_08998_)
  );
  sg13g2_o21ai_1 _18633_ (
    .A1(_08986_),
    .A2(_08988_),
    .B1(_08998_),
    .Y(_08999_)
  );
  sg13g2_nand2_1 _18634_ (
    .A(addr_i_4_),
    .B(_08266_),
    .Y(_09000_)
  );
  sg13g2_a22oi_1 _18635_ (
    .A1(_00159_),
    .A2(_09000_),
    .B1(_04276_),
    .B2(_00214_),
    .Y(_09001_)
  );
  sg13g2_nand2_1 _18636_ (
    .A(_00185_),
    .B(_02156_),
    .Y(_09002_)
  );
  sg13g2_nand2_1 _18637_ (
    .A(addr_i_3_),
    .B(_09002_),
    .Y(_09003_)
  );
  sg13g2_a21oi_1 _18638_ (
    .A1(addr_i_3_),
    .A2(_00194_),
    .B1(_09473_),
    .Y(_09004_)
  );
  sg13g2_nand2b_1 _18639_ (
    .A_N(_09004_),
    .B(addr_i_2_),
    .Y(_09005_)
  );
  sg13g2_a21oi_1 _18640_ (
    .A1(_00151_),
    .A2(_00926_),
    .B1(addr_i_3_),
    .Y(_09007_)
  );
  sg13g2_o21ai_1 _18641_ (
    .A1(_02330_),
    .A2(_09007_),
    .B1(_01279_),
    .Y(_09008_)
  );
  sg13g2_nand4_1 _18642_ (
    .A(_09001_),
    .B(_09003_),
    .C(_09005_),
    .D(_09008_),
    .Y(_09009_)
  );
  sg13g2_nand2_1 _18643_ (
    .A(_00744_),
    .B(_02349_),
    .Y(_09010_)
  );
  sg13g2_nand3_1 _18644_ (
    .A(addr_i_4_),
    .B(_00914_),
    .C(_01738_),
    .Y(_09011_)
  );
  sg13g2_o21ai_1 _18645_ (
    .A1(_06535_),
    .A2(_09010_),
    .B1(_09011_),
    .Y(_09012_)
  );
  sg13g2_a21oi_1 _18646_ (
    .A1(_00716_),
    .A2(_00975_),
    .B1(addr_i_3_),
    .Y(_09013_)
  );
  sg13g2_o21ai_1 _18647_ (
    .A1(_01972_),
    .A2(_09013_),
    .B1(addr_i_6_),
    .Y(_09014_)
  );
  sg13g2_o21ai_1 _18648_ (
    .A1(addr_i_6_),
    .A2(_09012_),
    .B1(_09014_),
    .Y(_09015_)
  );
  sg13g2_nor2_1 _18649_ (
    .A(_01041_),
    .B(_02443_),
    .Y(_09016_)
  );
  sg13g2_a21oi_1 _18650_ (
    .A1(_00148_),
    .A2(_01912_),
    .B1(addr_i_7_),
    .Y(_09018_)
  );
  sg13g2_o21ai_1 _18651_ (
    .A1(_03070_),
    .A2(_09018_),
    .B1(addr_i_3_),
    .Y(_09019_)
  );
  sg13g2_o21ai_1 _18652_ (
    .A1(addr_i_7_),
    .A2(_09016_),
    .B1(_09019_),
    .Y(_09020_)
  );
  sg13g2_o21ai_1 _18653_ (
    .A1(_09015_),
    .A2(_09020_),
    .B1(_02604_),
    .Y(_09021_)
  );
  sg13g2_and2_1 _18654_ (
    .A(_09009_),
    .B(_09021_),
    .X(_09022_)
  );
  sg13g2_a21oi_1 _18655_ (
    .A1(_08999_),
    .A2(_09022_),
    .B1(addr_i_10_),
    .Y(_09023_)
  );
  sg13g2_o21ai_1 _18656_ (
    .A1(_08976_),
    .A2(_09023_),
    .B1(_02251_),
    .Y(_09024_)
  );
  sg13g2_a21oi_1 _18657_ (
    .A1(addr_i_4_),
    .A2(_02405_),
    .B1(_05833_),
    .Y(_09025_)
  );
  sg13g2_nor2_1 _18658_ (
    .A(_03930_),
    .B(_09025_),
    .Y(_09026_)
  );
  sg13g2_a21oi_1 _18659_ (
    .A1(_01199_),
    .A2(_01499_),
    .B1(addr_i_4_),
    .Y(_09027_)
  );
  sg13g2_a22oi_1 _18660_ (
    .A1(_01365_),
    .A2(_00898_),
    .B1(_09026_),
    .B2(_09027_),
    .Y(_09028_)
  );
  sg13g2_nand2_1 _18661_ (
    .A(_02577_),
    .B(_00414_),
    .Y(_09029_)
  );
  sg13g2_a22oi_1 _18662_ (
    .A1(addr_i_4_),
    .A2(_09029_),
    .B1(_02014_),
    .B2(_00061_),
    .Y(_09030_)
  );
  sg13g2_a21o_1 _18663_ (
    .A1(_00048_),
    .A2(_09028_),
    .B1(_09030_),
    .X(_09031_)
  );
  sg13g2_nand2_1 _18664_ (
    .A(_00105_),
    .B(_01073_),
    .Y(_09032_)
  );
  sg13g2_a22oi_1 _18665_ (
    .A1(_06740_),
    .A2(_09032_),
    .B1(_05765_),
    .B2(addr_i_8_),
    .Y(_09033_)
  );
  sg13g2_o21ai_1 _18666_ (
    .A1(_01262_),
    .A2(_03690_),
    .B1(addr_i_3_),
    .Y(_09034_)
  );
  sg13g2_o21ai_1 _18667_ (
    .A1(addr_i_2_),
    .A2(_02448_),
    .B1(_09034_),
    .Y(_09035_)
  );
  sg13g2_o21ai_1 _18668_ (
    .A1(_04068_),
    .A2(_00561_),
    .B1(_06895_),
    .Y(_09036_)
  );
  sg13g2_o21ai_1 _18669_ (
    .A1(_02238_),
    .A2(_02976_),
    .B1(addr_i_3_),
    .Y(_09037_)
  );
  sg13g2_a21oi_1 _18670_ (
    .A1(_00764_),
    .A2(_09037_),
    .B1(addr_i_6_),
    .Y(_09040_)
  );
  sg13g2_a22oi_1 _18671_ (
    .A1(_01336_),
    .A2(_09036_),
    .B1(_09040_),
    .B2(_00257_),
    .Y(_09041_)
  );
  sg13g2_a21oi_1 _18672_ (
    .A1(addr_i_2_),
    .A2(_04246_),
    .B1(_02154_),
    .Y(_09042_)
  );
  sg13g2_nor2_1 _18673_ (
    .A(addr_i_3_),
    .B(_09042_),
    .Y(_09043_)
  );
  sg13g2_a22oi_1 _18674_ (
    .A1(_01191_),
    .A2(_00542_),
    .B1(_09043_),
    .B2(addr_i_4_),
    .Y(_09044_)
  );
  sg13g2_a21oi_1 _18675_ (
    .A1(addr_i_4_),
    .A2(_09041_),
    .B1(_09044_),
    .Y(_09045_)
  );
  sg13g2_a22oi_1 _18676_ (
    .A1(addr_i_6_),
    .A2(_09035_),
    .B1(_09045_),
    .B2(_00114_),
    .Y(_09046_)
  );
  sg13g2_a22oi_1 _18677_ (
    .A1(_09031_),
    .A2(_09033_),
    .B1(_00109_),
    .B2(_09046_),
    .Y(_09047_)
  );
  sg13g2_o21ai_1 _18678_ (
    .A1(_05645_),
    .A2(_04464_),
    .B1(addr_i_4_),
    .Y(_09048_)
  );
  sg13g2_a21oi_1 _18679_ (
    .A1(_01658_),
    .A2(_00353_),
    .B1(addr_i_4_),
    .Y(_09049_)
  );
  sg13g2_a22oi_1 _18680_ (
    .A1(addr_i_2_),
    .A2(_09002_),
    .B1(_09049_),
    .B2(_00301_),
    .Y(_09051_)
  );
  sg13g2_nand3_1 _18681_ (
    .A(addr_i_3_),
    .B(_09048_),
    .C(_09051_),
    .Y(_09052_)
  );
  sg13g2_o21ai_1 _18682_ (
    .A1(_02238_),
    .A2(_01542_),
    .B1(addr_i_4_),
    .Y(_09053_)
  );
  sg13g2_o21ai_1 _18683_ (
    .A1(addr_i_4_),
    .A2(_00911_),
    .B1(_09053_),
    .Y(_09054_)
  );
  sg13g2_or3_1 _18684_ (
    .A(addr_i_3_),
    .B(_07171_),
    .C(_09054_),
    .X(_09055_)
  );
  sg13g2_a22oi_1 _18685_ (
    .A1(_09052_),
    .A2(_09055_),
    .B1(_02040_),
    .B2(_01064_),
    .Y(_09056_)
  );
  sg13g2_a21o_1 _18686_ (
    .A1(addr_i_4_),
    .A2(_01949_),
    .B1(_03690_),
    .X(_09057_)
  );
  sg13g2_a21oi_1 _18687_ (
    .A1(addr_i_2_),
    .A2(_09057_),
    .B1(_09027_),
    .Y(_09058_)
  );
  sg13g2_o21ai_1 _18688_ (
    .A1(addr_i_5_),
    .A2(_06927_),
    .B1(_01450_),
    .Y(_09059_)
  );
  sg13g2_nand3_1 _18689_ (
    .A(_00056_),
    .B(_02822_),
    .C(_09059_),
    .Y(_09060_)
  );
  sg13g2_o21ai_1 _18690_ (
    .A1(_00105_),
    .A2(_00402_),
    .B1(_08492_),
    .Y(_09062_)
  );
  sg13g2_a221oi_1 _18691_ (
    .A1(addr_i_2_),
    .A2(_09060_),
    .B1(_09062_),
    .B2(_00239_),
    .C1(_04036_),
    .Y(_09063_)
  );
  sg13g2_o21ai_1 _18692_ (
    .A1(addr_i_3_),
    .A2(_09058_),
    .B1(_09063_),
    .Y(_09064_)
  );
  sg13g2_nand2_1 _18693_ (
    .A(addr_i_11_),
    .B(_09064_),
    .Y(_09065_)
  );
  sg13g2_o21ai_1 _18694_ (
    .A1(_01308_),
    .A2(_04367_),
    .B1(_01524_),
    .Y(_09066_)
  );
  sg13g2_a221oi_1 _18695_ (
    .A1(addr_i_3_),
    .A2(_05769_),
    .B1(_09066_),
    .B2(addr_i_7_),
    .C1(_01064_),
    .Y(_09067_)
  );
  sg13g2_a21oi_1 _18696_ (
    .A1(_07458_),
    .A2(_02200_),
    .B1(_06518_),
    .Y(_09068_)
  );
  sg13g2_nand2_1 _18697_ (
    .A(_07284_),
    .B(_09068_),
    .Y(_09069_)
  );
  sg13g2_o21ai_1 _18698_ (
    .A1(addr_i_3_),
    .A2(_00118_),
    .B1(_00573_),
    .Y(_09070_)
  );
  sg13g2_a221oi_1 _18699_ (
    .A1(addr_i_5_),
    .A2(_09069_),
    .B1(_09070_),
    .B2(_00292_),
    .C1(_01819_),
    .Y(_09071_)
  );
  sg13g2_o21ai_1 _18700_ (
    .A1(addr_i_4_),
    .A2(_09067_),
    .B1(_09071_),
    .Y(_09073_)
  );
  sg13g2_a21oi_1 _18701_ (
    .A1(_00414_),
    .A2(_04799_),
    .B1(addr_i_3_),
    .Y(_09074_)
  );
  sg13g2_a21oi_1 _18702_ (
    .A1(_07724_),
    .A2(_01224_),
    .B1(addr_i_2_),
    .Y(_09075_)
  );
  sg13g2_nor3_1 _18703_ (
    .A(_06010_),
    .B(_00315_),
    .C(_00206_),
    .Y(_09076_)
  );
  sg13g2_nor4_1 _18704_ (
    .A(_00802_),
    .B(_09074_),
    .C(_09075_),
    .D(_09076_),
    .Y(_09077_)
  );
  sg13g2_a21o_1 _18705_ (
    .A1(addr_i_2_),
    .A2(_01765_),
    .B1(_00128_),
    .X(_09078_)
  );
  sg13g2_a21oi_1 _18706_ (
    .A1(_02528_),
    .A2(_00820_),
    .B1(_01520_),
    .Y(_09079_)
  );
  sg13g2_a21oi_1 _18707_ (
    .A1(_05877_),
    .A2(_09078_),
    .B1(_09079_),
    .Y(_09080_)
  );
  sg13g2_and2_1 _18708_ (
    .A(_01131_),
    .B(_03637_),
    .X(_09081_)
  );
  sg13g2_o21ai_1 _18709_ (
    .A1(_00617_),
    .A2(_09081_),
    .B1(addr_i_3_),
    .Y(_09082_)
  );
  sg13g2_a21oi_1 _18710_ (
    .A1(_09080_),
    .A2(_09082_),
    .B1(_01082_),
    .Y(_09084_)
  );
  sg13g2_a22oi_1 _18711_ (
    .A1(addr_i_8_),
    .A2(_09073_),
    .B1(_09077_),
    .B2(_09084_),
    .Y(_09085_)
  );
  sg13g2_a21oi_1 _18712_ (
    .A1(_08752_),
    .A2(_02405_),
    .B1(_01191_),
    .Y(_09086_)
  );
  sg13g2_o21ai_1 _18713_ (
    .A1(addr_i_4_),
    .A2(_09086_),
    .B1(_04534_),
    .Y(_09087_)
  );
  sg13g2_nor2_1 _18714_ (
    .A(_05218_),
    .B(_01957_),
    .Y(_09088_)
  );
  sg13g2_nand2_1 _18715_ (
    .A(_01353_),
    .B(_07724_),
    .Y(_09089_)
  );
  sg13g2_a22oi_1 _18716_ (
    .A1(addr_i_3_),
    .A2(_09089_),
    .B1(_02391_),
    .B2(addr_i_7_),
    .Y(_09090_)
  );
  sg13g2_a21oi_1 _18717_ (
    .A1(_00916_),
    .A2(_09088_),
    .B1(_09090_),
    .Y(_09091_)
  );
  sg13g2_a22oi_1 _18718_ (
    .A1(_00068_),
    .A2(_09087_),
    .B1(_09091_),
    .B2(_01151_),
    .Y(_09092_)
  );
  sg13g2_nand2_1 _18719_ (
    .A(addr_i_3_),
    .B(_07871_),
    .Y(_09093_)
  );
  sg13g2_nand3_1 _18720_ (
    .A(_02930_),
    .B(_00077_),
    .C(_09093_),
    .Y(_09095_)
  );
  sg13g2_nor3_1 _18721_ (
    .A(_00065_),
    .B(addr_i_5_),
    .C(_01086_),
    .Y(_09096_)
  );
  sg13g2_a22oi_1 _18722_ (
    .A1(addr_i_3_),
    .A2(_00080_),
    .B1(_09096_),
    .B2(addr_i_7_),
    .Y(_09097_)
  );
  sg13g2_nor3_1 _18723_ (
    .A(_04068_),
    .B(_02203_),
    .C(_02935_),
    .Y(_09098_)
  );
  sg13g2_o21ai_1 _18724_ (
    .A1(addr_i_2_),
    .A2(_00607_),
    .B1(_00838_),
    .Y(_09099_)
  );
  sg13g2_o21ai_1 _18725_ (
    .A1(_09097_),
    .A2(_09098_),
    .B1(_09099_),
    .Y(_09100_)
  );
  sg13g2_a22oi_1 _18726_ (
    .A1(addr_i_5_),
    .A2(_09095_),
    .B1(_09100_),
    .B2(addr_i_8_),
    .Y(_09101_)
  );
  sg13g2_nor2_1 _18727_ (
    .A(_09092_),
    .B(_09101_),
    .Y(_09102_)
  );
  sg13g2_nor2_1 _18728_ (
    .A(addr_i_9_),
    .B(_09102_),
    .Y(_09103_)
  );
  sg13g2_a22oi_1 _18729_ (
    .A1(addr_i_9_),
    .A2(_09085_),
    .B1(_09103_),
    .B2(addr_i_10_),
    .Y(_09104_)
  );
  sg13g2_nor4_1 _18730_ (
    .A(_09047_),
    .B(_09056_),
    .C(_09065_),
    .D(_09104_),
    .Y(_09106_)
  );
  sg13g2_o21ai_1 _18731_ (
    .A1(_01616_),
    .A2(_01127_),
    .B1(_04442_),
    .Y(_09107_)
  );
  sg13g2_a21oi_1 _18732_ (
    .A1(_01473_),
    .A2(_02887_),
    .B1(_00951_),
    .Y(_09108_)
  );
  sg13g2_o21ai_1 _18733_ (
    .A1(_01580_),
    .A2(_09108_),
    .B1(addr_i_2_),
    .Y(_09109_)
  );
  sg13g2_nand2_1 _18734_ (
    .A(_00483_),
    .B(_00759_),
    .Y(_09110_)
  );
  sg13g2_a21oi_1 _18735_ (
    .A1(_01843_),
    .A2(_09110_),
    .B1(_08388_),
    .Y(_09111_)
  );
  sg13g2_o21ai_1 _18736_ (
    .A1(addr_i_7_),
    .A2(_01244_),
    .B1(_00744_),
    .Y(_09112_)
  );
  sg13g2_nand2_1 _18737_ (
    .A(_03358_),
    .B(_09112_),
    .Y(_09113_)
  );
  sg13g2_o21ai_1 _18738_ (
    .A1(_09111_),
    .A2(_09113_),
    .B1(_02796_),
    .Y(_09114_)
  );
  sg13g2_nand4_1 _18739_ (
    .A(_01692_),
    .B(_09107_),
    .C(_09109_),
    .D(_09114_),
    .Y(_09115_)
  );
  sg13g2_o21ai_1 _18740_ (
    .A1(_02976_),
    .A2(_01604_),
    .B1(addr_i_3_),
    .Y(_09117_)
  );
  sg13g2_nand3_1 _18741_ (
    .A(_00994_),
    .B(_02694_),
    .C(_09117_),
    .Y(_09118_)
  );
  sg13g2_a21oi_1 _18742_ (
    .A1(addr_i_3_),
    .A2(_09448_),
    .B1(_01091_),
    .Y(_09119_)
  );
  sg13g2_o21ai_1 _18743_ (
    .A1(addr_i_7_),
    .A2(_09119_),
    .B1(_00629_),
    .Y(_09120_)
  );
  sg13g2_a21oi_1 _18744_ (
    .A1(addr_i_2_),
    .A2(_01588_),
    .B1(_00445_),
    .Y(_09121_)
  );
  sg13g2_nor2_1 _18745_ (
    .A(_00838_),
    .B(_09121_),
    .Y(_09122_)
  );
  sg13g2_nor3_1 _18746_ (
    .A(addr_i_7_),
    .B(_06806_),
    .C(_00399_),
    .Y(_09123_)
  );
  sg13g2_a22oi_1 _18747_ (
    .A1(addr_i_7_),
    .A2(_09122_),
    .B1(_09123_),
    .B2(addr_i_3_),
    .Y(_09124_)
  );
  sg13g2_a22oi_1 _18748_ (
    .A1(_01630_),
    .A2(_09118_),
    .B1(_09120_),
    .B2(_09124_),
    .Y(_09125_)
  );
  sg13g2_a21oi_1 _18749_ (
    .A1(addr_i_8_),
    .A2(_09115_),
    .B1(_09125_),
    .Y(_09126_)
  );
  sg13g2_o21ai_1 _18750_ (
    .A1(addr_i_2_),
    .A2(_08930_),
    .B1(_02832_),
    .Y(_09128_)
  );
  sg13g2_a21oi_1 _18751_ (
    .A1(_00380_),
    .A2(_01273_),
    .B1(addr_i_3_),
    .Y(_09129_)
  );
  sg13g2_a22oi_1 _18752_ (
    .A1(addr_i_4_),
    .A2(_09128_),
    .B1(_09129_),
    .B2(_00206_),
    .Y(_09130_)
  );
  sg13g2_nand3_1 _18753_ (
    .A(addr_i_7_),
    .B(_07610_),
    .C(_09130_),
    .Y(_09131_)
  );
  sg13g2_a21oi_1 _18754_ (
    .A1(_00155_),
    .A2(_08020_),
    .B1(addr_i_4_),
    .Y(_09132_)
  );
  sg13g2_or2_1 _18755_ (
    .A(_09348_),
    .B(_09129_),
    .X(_09133_)
  );
  sg13g2_o21ai_1 _18756_ (
    .A1(_09132_),
    .A2(_09133_),
    .B1(_01475_),
    .Y(_09134_)
  );
  sg13g2_nand3_1 _18757_ (
    .A(addr_i_8_),
    .B(_09131_),
    .C(_09134_),
    .Y(_09135_)
  );
  sg13g2_o21ai_1 _18758_ (
    .A1(addr_i_3_),
    .A2(_01972_),
    .B1(_09492_),
    .Y(_09136_)
  );
  sg13g2_a21oi_1 _18759_ (
    .A1(_00930_),
    .A2(_00688_),
    .B1(_00485_),
    .Y(_09137_)
  );
  sg13g2_a221oi_1 _18760_ (
    .A1(_01262_),
    .A2(_00298_),
    .B1(_09136_),
    .B2(_04191_),
    .C1(_09137_),
    .Y(_09139_)
  );
  sg13g2_nor4_1 _18761_ (
    .A(addr_i_7_),
    .B(_01459_),
    .C(_00960_),
    .D(_06804_),
    .Y(_09140_)
  );
  sg13g2_o21ai_1 _18762_ (
    .A1(_01472_),
    .A2(_06176_),
    .B1(_02387_),
    .Y(_09141_)
  );
  sg13g2_a21oi_1 _18763_ (
    .A1(_01029_),
    .A2(_09141_),
    .B1(_08708_),
    .Y(_09142_)
  );
  sg13g2_nand2_1 _18764_ (
    .A(addr_i_3_),
    .B(_00183_),
    .Y(_09143_)
  );
  sg13g2_a21oi_1 _18765_ (
    .A1(_01008_),
    .A2(_09143_),
    .B1(_03431_),
    .Y(_09144_)
  );
  sg13g2_nor4_1 _18766_ (
    .A(addr_i_8_),
    .B(_09140_),
    .C(_09142_),
    .D(_09144_),
    .Y(_09145_)
  );
  sg13g2_o21ai_1 _18767_ (
    .A1(_02257_),
    .A2(_09139_),
    .B1(_09145_),
    .Y(_09146_)
  );
  sg13g2_nand3_1 _18768_ (
    .A(addr_i_9_),
    .B(_09135_),
    .C(_09146_),
    .Y(_09147_)
  );
  sg13g2_o21ai_1 _18769_ (
    .A1(addr_i_9_),
    .A2(_09126_),
    .B1(_09147_),
    .Y(_09148_)
  );
  sg13g2_nor2_1 _18770_ (
    .A(addr_i_10_),
    .B(_09148_),
    .Y(_09151_)
  );
  sg13g2_a22oi_1 _18771_ (
    .A1(_09105_),
    .A2(_02380_),
    .B1(_02179_),
    .B2(_03073_),
    .Y(_09152_)
  );
  sg13g2_a22oi_1 _18772_ (
    .A1(_00403_),
    .A2(_00315_),
    .B1(_01191_),
    .B2(_01630_),
    .Y(_09153_)
  );
  sg13g2_a21oi_1 _18773_ (
    .A1(_01630_),
    .A2(_06536_),
    .B1(_09153_),
    .Y(_09154_)
  );
  sg13g2_a21oi_1 _18774_ (
    .A1(_00391_),
    .A2(_01499_),
    .B1(addr_i_3_),
    .Y(_09155_)
  );
  sg13g2_a21oi_1 _18775_ (
    .A1(_00077_),
    .A2(_00470_),
    .B1(addr_i_2_),
    .Y(_09156_)
  );
  sg13g2_nor4_1 _18776_ (
    .A(_07171_),
    .B(_04036_),
    .C(_09155_),
    .D(_09156_),
    .Y(_09157_)
  );
  sg13g2_a221oi_1 _18777_ (
    .A1(_05313_),
    .A2(_09152_),
    .B1(_09154_),
    .B2(_09157_),
    .C1(addr_i_11_),
    .Y(_09158_)
  );
  sg13g2_nand3_1 _18778_ (
    .A(addr_i_5_),
    .B(_01367_),
    .C(_06070_),
    .Y(_09159_)
  );
  sg13g2_nor2_1 _18779_ (
    .A(_05877_),
    .B(_04139_),
    .Y(_09160_)
  );
  sg13g2_a22oi_1 _18780_ (
    .A1(addr_i_6_),
    .A2(_03839_),
    .B1(_01869_),
    .B2(addr_i_3_),
    .Y(_09162_)
  );
  sg13g2_a22oi_1 _18781_ (
    .A1(_09159_),
    .A2(_09160_),
    .B1(_09162_),
    .B2(addr_i_7_),
    .Y(_09163_)
  );
  sg13g2_a22oi_1 _18782_ (
    .A1(addr_i_3_),
    .A2(_02304_),
    .B1(_00279_),
    .B2(_07889_),
    .Y(_09164_)
  );
  sg13g2_nand2b_1 _18783_ (
    .A_N(_09164_),
    .B(addr_i_7_),
    .Y(_09165_)
  );
  sg13g2_a21oi_1 _18784_ (
    .A1(_05479_),
    .A2(_09165_),
    .B1(addr_i_6_),
    .Y(_09166_)
  );
  sg13g2_o21ai_1 _18785_ (
    .A1(_09163_),
    .A2(_09166_),
    .B1(_01350_),
    .Y(_09167_)
  );
  sg13g2_nor3_1 _18786_ (
    .A(_00053_),
    .B(_03308_),
    .C(_04939_),
    .Y(_09168_)
  );
  sg13g2_o21ai_1 _18787_ (
    .A1(_07824_),
    .A2(_00815_),
    .B1(_00544_),
    .Y(_09169_)
  );
  sg13g2_nor2_1 _18788_ (
    .A(_02089_),
    .B(_05805_),
    .Y(_09170_)
  );
  sg13g2_a22oi_1 _18789_ (
    .A1(_01892_),
    .A2(_09169_),
    .B1(_09170_),
    .B2(_07293_),
    .Y(_09171_)
  );
  sg13g2_a21oi_1 _18790_ (
    .A1(_02297_),
    .A2(_00884_),
    .B1(_04052_),
    .Y(_09173_)
  );
  sg13g2_o21ai_1 _18791_ (
    .A1(_05266_),
    .A2(_09173_),
    .B1(_06630_),
    .Y(_09174_)
  );
  sg13g2_nand2_1 _18792_ (
    .A(_09171_),
    .B(_09174_),
    .Y(_09175_)
  );
  sg13g2_nor2_1 _18793_ (
    .A(addr_i_2_),
    .B(_03348_),
    .Y(_09176_)
  );
  sg13g2_o21ai_1 _18794_ (
    .A1(addr_i_4_),
    .A2(_09176_),
    .B1(_00504_),
    .Y(_09177_)
  );
  sg13g2_nand3_1 _18795_ (
    .A(addr_i_3_),
    .B(addr_i_5_),
    .C(_00408_),
    .Y(_09178_)
  );
  sg13g2_o21ai_1 _18796_ (
    .A1(addr_i_3_),
    .A2(_00815_),
    .B1(_09178_),
    .Y(_09179_)
  );
  sg13g2_a221oi_1 _18797_ (
    .A1(_00529_),
    .A2(_09177_),
    .B1(_09179_),
    .B2(_09138_),
    .C1(addr_i_8_),
    .Y(_09180_)
  );
  sg13g2_a21o_1 _18798_ (
    .A1(addr_i_4_),
    .A2(_03485_),
    .B1(_00644_),
    .X(_09181_)
  );
  sg13g2_o21ai_1 _18799_ (
    .A1(_03267_),
    .A2(_01376_),
    .B1(addr_i_6_),
    .Y(_09182_)
  );
  sg13g2_nand2b_1 _18800_ (
    .A_N(_09181_),
    .B(_09182_),
    .Y(_09184_)
  );
  sg13g2_nand2_1 _18801_ (
    .A(_06630_),
    .B(_09184_),
    .Y(_09185_)
  );
  sg13g2_a21oi_1 _18802_ (
    .A1(_09180_),
    .A2(_09185_),
    .B1(_00925_),
    .Y(_09186_)
  );
  sg13g2_o21ai_1 _18803_ (
    .A1(_09168_),
    .A2(_09175_),
    .B1(_09186_),
    .Y(_09187_)
  );
  sg13g2_nand3_1 _18804_ (
    .A(_09158_),
    .B(_09167_),
    .C(_09187_),
    .Y(_09188_)
  );
  sg13g2_nand2_1 _18805_ (
    .A(_02268_),
    .B(_04426_),
    .Y(_09189_)
  );
  sg13g2_o21ai_1 _18806_ (
    .A1(_00403_),
    .A2(_07643_),
    .B1(_09189_),
    .Y(_09190_)
  );
  sg13g2_nor3_1 _18807_ (
    .A(_04672_),
    .B(_01025_),
    .C(_04130_),
    .Y(_09191_)
  );
  sg13g2_a21oi_1 _18808_ (
    .A1(_08084_),
    .A2(_03428_),
    .B1(_02179_),
    .Y(_09192_)
  );
  sg13g2_a22oi_1 _18809_ (
    .A1(addr_i_4_),
    .A2(_01861_),
    .B1(_09192_),
    .B2(addr_i_9_),
    .Y(_09193_)
  );
  sg13g2_nand2_1 _18810_ (
    .A(_00697_),
    .B(_00080_),
    .Y(_09195_)
  );
  sg13g2_nand3_1 _18811_ (
    .A(addr_i_3_),
    .B(addr_i_6_),
    .C(_06032_),
    .Y(_09196_)
  );
  sg13g2_a21oi_1 _18812_ (
    .A1(_07706_),
    .A2(_09196_),
    .B1(_08708_),
    .Y(_09197_)
  );
  sg13g2_a22oi_1 _18813_ (
    .A1(_00128_),
    .A2(_09195_),
    .B1(_09197_),
    .B2(_07403_),
    .Y(_09198_)
  );
  sg13g2_o21ai_1 _18814_ (
    .A1(addr_i_5_),
    .A2(_02536_),
    .B1(_03871_),
    .Y(_09199_)
  );
  sg13g2_a21oi_1 _18815_ (
    .A1(_00388_),
    .A2(_09199_),
    .B1(_07614_),
    .Y(_09200_)
  );
  sg13g2_nor2_1 _18816_ (
    .A(_09198_),
    .B(_09200_),
    .Y(_09201_)
  );
  sg13g2_nand3b_1 _18817_ (
    .A_N(_09191_),
    .B(_09193_),
    .C(_09201_),
    .Y(_09202_)
  );
  sg13g2_a21oi_1 _18818_ (
    .A1(addr_i_9_),
    .A2(_02397_),
    .B1(addr_i_10_),
    .Y(_09203_)
  );
  sg13g2_a221oi_1 _18819_ (
    .A1(_03084_),
    .A2(_09190_),
    .B1(_09202_),
    .B2(_09203_),
    .C1(_01640_),
    .Y(_09204_)
  );
  sg13g2_nor2_1 _18820_ (
    .A(_00812_),
    .B(_09204_),
    .Y(_09206_)
  );
  sg13g2_o21ai_1 _18821_ (
    .A1(_09151_),
    .A2(_09188_),
    .B1(_09206_),
    .Y(_09207_)
  );
  sg13g2_o21ai_1 _18822_ (
    .A1(_09024_),
    .A2(_09106_),
    .B1(_09207_),
    .Y(data_o_8_)
  );
  sg13g2_o21ai_1 _18823_ (
    .A1(addr_i_6_),
    .A2(_00386_),
    .B1(_00122_),
    .Y(_09208_)
  );
  sg13g2_nand3_1 _18824_ (
    .A(addr_i_5_),
    .B(_00825_),
    .C(_09208_),
    .Y(_09209_)
  );
  sg13g2_or3_1 _18825_ (
    .A(addr_i_5_),
    .B(_00096_),
    .C(_07947_),
    .X(_09210_)
  );
  sg13g2_nand3_1 _18826_ (
    .A(_00061_),
    .B(_09209_),
    .C(_09210_),
    .Y(_09211_)
  );
  sg13g2_nand2_1 _18827_ (
    .A(_00616_),
    .B(_06223_),
    .Y(_09212_)
  );
  sg13g2_nand3_1 _18828_ (
    .A(_08232_),
    .B(_01411_),
    .C(_09212_),
    .Y(_09213_)
  );
  sg13g2_a21oi_1 _18829_ (
    .A1(_06784_),
    .A2(_00405_),
    .B1(_02191_),
    .Y(_09214_)
  );
  sg13g2_a22oi_1 _18830_ (
    .A1(addr_i_4_),
    .A2(_09213_),
    .B1(_09214_),
    .B2(addr_i_8_),
    .Y(_09216_)
  );
  sg13g2_nand3_1 _18831_ (
    .A(addr_i_6_),
    .B(_03424_),
    .C(_03853_),
    .Y(_09217_)
  );
  sg13g2_o21ai_1 _18832_ (
    .A1(_00840_),
    .A2(_00898_),
    .B1(addr_i_4_),
    .Y(_09218_)
  );
  sg13g2_nand2_1 _18833_ (
    .A(_09217_),
    .B(_09218_),
    .Y(_09219_)
  );
  sg13g2_o21ai_1 _18834_ (
    .A1(_00230_),
    .A2(_02304_),
    .B1(addr_i_8_),
    .Y(_09220_)
  );
  sg13g2_nand2_1 _18835_ (
    .A(addr_i_7_),
    .B(_08520_),
    .Y(_09221_)
  );
  sg13g2_nor2_1 _18836_ (
    .A(addr_i_2_),
    .B(_09221_),
    .Y(_09222_)
  );
  sg13g2_nand3_1 _18837_ (
    .A(_00200_),
    .B(_01008_),
    .C(_01343_),
    .Y(_09223_)
  );
  sg13g2_o21ai_1 _18838_ (
    .A1(_00074_),
    .A2(_09222_),
    .B1(_09223_),
    .Y(_09224_)
  );
  sg13g2_nand2_1 _18839_ (
    .A(addr_i_4_),
    .B(_08977_),
    .Y(_09225_)
  );
  sg13g2_a21oi_1 _18840_ (
    .A1(_09224_),
    .A2(_09225_),
    .B1(_00116_),
    .Y(_09227_)
  );
  sg13g2_a22oi_1 _18841_ (
    .A1(_00061_),
    .A2(_09219_),
    .B1(_09220_),
    .B2(_09227_),
    .Y(_09228_)
  );
  sg13g2_a22oi_1 _18842_ (
    .A1(_09211_),
    .A2(_09216_),
    .B1(_09326_),
    .B2(_09228_),
    .Y(_09229_)
  );
  sg13g2_nor2_1 _18843_ (
    .A(addr_i_7_),
    .B(_03737_),
    .Y(_09230_)
  );
  sg13g2_a221oi_1 _18844_ (
    .A1(_06927_),
    .A2(_08180_),
    .B1(_03766_),
    .B2(_00183_),
    .C1(_09230_),
    .Y(_09231_)
  );
  sg13g2_nand2_1 _18845_ (
    .A(_01672_),
    .B(_07359_),
    .Y(_09232_)
  );
  sg13g2_o21ai_1 _18846_ (
    .A1(_00959_),
    .A2(_06132_),
    .B1(_09232_),
    .Y(_09233_)
  );
  sg13g2_a221oi_1 _18847_ (
    .A1(_01191_),
    .A2(_01998_),
    .B1(_09233_),
    .B2(_00949_),
    .C1(addr_i_3_),
    .Y(_09234_)
  );
  sg13g2_a21o_1 _18848_ (
    .A1(addr_i_3_),
    .A2(_09231_),
    .B1(_09234_),
    .X(_09235_)
  );
  sg13g2_o21ai_1 _18849_ (
    .A1(_04307_),
    .A2(_04082_),
    .B1(_02271_),
    .Y(_09236_)
  );
  sg13g2_nand3_1 _18850_ (
    .A(addr_i_3_),
    .B(addr_i_7_),
    .C(_03452_),
    .Y(_09238_)
  );
  sg13g2_nand2_1 _18851_ (
    .A(_09236_),
    .B(_09238_),
    .Y(_09239_)
  );
  sg13g2_o21ai_1 _18852_ (
    .A1(_00792_),
    .A2(_01016_),
    .B1(addr_i_5_),
    .Y(_09240_)
  );
  sg13g2_o21ai_1 _18853_ (
    .A1(_04068_),
    .A2(_08598_),
    .B1(_00561_),
    .Y(_09241_)
  );
  sg13g2_o21ai_1 _18854_ (
    .A1(_00536_),
    .A2(_01551_),
    .B1(_00305_),
    .Y(_09242_)
  );
  sg13g2_nand4_1 _18855_ (
    .A(_00113_),
    .B(_09240_),
    .C(_09241_),
    .D(_09242_),
    .Y(_09243_)
  );
  sg13g2_a21oi_1 _18856_ (
    .A1(addr_i_6_),
    .A2(_09239_),
    .B1(_09243_),
    .Y(_09244_)
  );
  sg13g2_a22oi_1 _18857_ (
    .A1(addr_i_8_),
    .A2(_09235_),
    .B1(_09244_),
    .B2(addr_i_9_),
    .Y(_09245_)
  );
  sg13g2_o21ai_1 _18858_ (
    .A1(_09229_),
    .A2(_09245_),
    .B1(_01774_),
    .Y(_09246_)
  );
  sg13g2_a21oi_1 _18859_ (
    .A1(_00561_),
    .A2(_00542_),
    .B1(_04555_),
    .Y(_09247_)
  );
  sg13g2_o21ai_1 _18860_ (
    .A1(addr_i_4_),
    .A2(_09247_),
    .B1(_08704_),
    .Y(_09249_)
  );
  sg13g2_a21o_1 _18861_ (
    .A1(_03669_),
    .A2(_07288_),
    .B1(_00067_),
    .X(_09250_)
  );
  sg13g2_nand3_1 _18862_ (
    .A(_02898_),
    .B(_03754_),
    .C(_00595_),
    .Y(_09251_)
  );
  sg13g2_a22oi_1 _18863_ (
    .A1(_04191_),
    .A2(_09251_),
    .B1(_00334_),
    .B2(_00351_),
    .Y(_09252_)
  );
  sg13g2_a21oi_1 _18864_ (
    .A1(_09250_),
    .A2(_09252_),
    .B1(_00367_),
    .Y(_09253_)
  );
  sg13g2_o21ai_1 _18865_ (
    .A1(addr_i_2_),
    .A2(_00412_),
    .B1(_00276_),
    .Y(_09254_)
  );
  sg13g2_a21oi_1 _18866_ (
    .A1(_00185_),
    .A2(_02497_),
    .B1(addr_i_3_),
    .Y(_09255_)
  );
  sg13g2_a22oi_1 _18867_ (
    .A1(addr_i_3_),
    .A2(_09181_),
    .B1(_09254_),
    .B2(_09255_),
    .Y(_09256_)
  );
  sg13g2_or4_1 _18868_ (
    .A(addr_i_6_),
    .B(_01445_),
    .C(_07603_),
    .D(_03188_),
    .X(_09257_)
  );
  sg13g2_nand3_1 _18869_ (
    .A(_00344_),
    .B(_01382_),
    .C(_02028_),
    .Y(_09258_)
  );
  sg13g2_nand3_1 _18870_ (
    .A(addr_i_9_),
    .B(_09257_),
    .C(_09258_),
    .Y(_09261_)
  );
  sg13g2_a22oi_1 _18871_ (
    .A1(_09249_),
    .A2(_09253_),
    .B1(_09256_),
    .B2(_09261_),
    .Y(_09262_)
  );
  sg13g2_nor2_1 _18872_ (
    .A(addr_i_3_),
    .B(_07744_),
    .Y(_09263_)
  );
  sg13g2_a21oi_1 _18873_ (
    .A1(addr_i_3_),
    .A2(_01543_),
    .B1(_09263_),
    .Y(_09264_)
  );
  sg13g2_a21oi_1 _18874_ (
    .A1(_00069_),
    .A2(_02810_),
    .B1(_09491_),
    .Y(_09265_)
  );
  sg13g2_a21oi_1 _18875_ (
    .A1(_09094_),
    .A2(_00645_),
    .B1(_09265_),
    .Y(_09266_)
  );
  sg13g2_o21ai_1 _18876_ (
    .A1(addr_i_2_),
    .A2(_09264_),
    .B1(_09266_),
    .Y(_09267_)
  );
  sg13g2_a21oi_1 _18877_ (
    .A1(_06779_),
    .A2(_03179_),
    .B1(addr_i_7_),
    .Y(_09268_)
  );
  sg13g2_a21oi_1 _18878_ (
    .A1(addr_i_6_),
    .A2(_09267_),
    .B1(_09268_),
    .Y(_09269_)
  );
  sg13g2_nand4_1 _18879_ (
    .A(addr_i_3_),
    .B(_00482_),
    .C(_00353_),
    .D(_02560_),
    .Y(_09270_)
  );
  sg13g2_a21oi_1 _18880_ (
    .A1(_05402_),
    .A2(_00591_),
    .B1(_08732_),
    .Y(_09272_)
  );
  sg13g2_nand2_1 _18881_ (
    .A(_00190_),
    .B(_09272_),
    .Y(_09273_)
  );
  sg13g2_a21oi_1 _18882_ (
    .A1(_09270_),
    .A2(_09273_),
    .B1(_08674_),
    .Y(_09274_)
  );
  sg13g2_nor2_1 _18883_ (
    .A(_00827_),
    .B(_00279_),
    .Y(_09275_)
  );
  sg13g2_a21oi_1 _18884_ (
    .A1(_00771_),
    .A2(_09275_),
    .B1(_04672_),
    .Y(_09276_)
  );
  sg13g2_o21ai_1 _18885_ (
    .A1(_00666_),
    .A2(_05544_),
    .B1(_01666_),
    .Y(_09277_)
  );
  sg13g2_a22oi_1 _18886_ (
    .A1(_02528_),
    .A2(_01227_),
    .B1(_00794_),
    .B2(_09277_),
    .Y(_09278_)
  );
  sg13g2_nor4_1 _18887_ (
    .A(addr_i_9_),
    .B(_09274_),
    .C(_09276_),
    .D(_09278_),
    .Y(_09279_)
  );
  sg13g2_o21ai_1 _18888_ (
    .A1(addr_i_8_),
    .A2(_09269_),
    .B1(_09279_),
    .Y(_09280_)
  );
  sg13g2_nand3b_1 _18889_ (
    .A_N(_09262_),
    .B(addr_i_10_),
    .C(_09280_),
    .Y(_09281_)
  );
  sg13g2_nand3_1 _18890_ (
    .A(_03051_),
    .B(_09246_),
    .C(_09281_),
    .Y(_09283_)
  );
  sg13g2_a221oi_1 _18891_ (
    .A1(_01282_),
    .A2(_00262_),
    .B1(_01508_),
    .B2(_00786_),
    .C1(_06361_),
    .Y(_09284_)
  );
  sg13g2_o21ai_1 _18892_ (
    .A1(_05252_),
    .A2(_07871_),
    .B1(addr_i_5_),
    .Y(_09285_)
  );
  sg13g2_and3_1 _18893_ (
    .A(addr_i_3_),
    .B(_04109_),
    .C(_09285_),
    .X(_09286_)
  );
  sg13g2_a21oi_1 _18894_ (
    .A1(_00061_),
    .A2(_09284_),
    .B1(_09286_),
    .Y(_09287_)
  );
  sg13g2_a21oi_1 _18895_ (
    .A1(_02513_),
    .A2(_01224_),
    .B1(addr_i_2_),
    .Y(_09288_)
  );
  sg13g2_o21ai_1 _18896_ (
    .A1(_03906_),
    .A2(_09288_),
    .B1(addr_i_3_),
    .Y(_09289_)
  );
  sg13g2_a22oi_1 _18897_ (
    .A1(_03150_),
    .A2(_03190_),
    .B1(_04062_),
    .B2(_00290_),
    .Y(_09290_)
  );
  sg13g2_a21oi_1 _18898_ (
    .A1(_09289_),
    .A2(_09290_),
    .B1(_02718_),
    .Y(_09291_)
  );
  sg13g2_o21ai_1 _18899_ (
    .A1(addr_i_8_),
    .A2(_09287_),
    .B1(_09291_),
    .Y(_09292_)
  );
  sg13g2_nor2_1 _18900_ (
    .A(addr_i_10_),
    .B(_05659_),
    .Y(_09294_)
  );
  sg13g2_a22oi_1 _18901_ (
    .A1(_00945_),
    .A2(_02578_),
    .B1(_02542_),
    .B2(_05834_),
    .Y(_09295_)
  );
  sg13g2_nor3_1 _18902_ (
    .A(_03690_),
    .B(_02040_),
    .C(_09295_),
    .Y(_09296_)
  );
  sg13g2_a22oi_1 _18903_ (
    .A1(_09292_),
    .A2(_09294_),
    .B1(_09296_),
    .B2(_01640_),
    .Y(_09297_)
  );
  sg13g2_nor2_1 _18904_ (
    .A(_00812_),
    .B(_09297_),
    .Y(_09298_)
  );
  sg13g2_nand3_1 _18905_ (
    .A(addr_i_4_),
    .B(_01290_),
    .C(_01709_),
    .Y(_09299_)
  );
  sg13g2_o21ai_1 _18906_ (
    .A1(addr_i_4_),
    .A2(_02008_),
    .B1(_09299_),
    .Y(_09300_)
  );
  sg13g2_nor2_1 _18907_ (
    .A(_08487_),
    .B(_03899_),
    .Y(_09301_)
  );
  sg13g2_o21ai_1 _18908_ (
    .A1(_01888_),
    .A2(_01014_),
    .B1(addr_i_3_),
    .Y(_09302_)
  );
  sg13g2_a21oi_1 _18909_ (
    .A1(_00224_),
    .A2(_09302_),
    .B1(addr_i_5_),
    .Y(_09303_)
  );
  sg13g2_a22oi_1 _18910_ (
    .A1(_07824_),
    .A2(_04747_),
    .B1(_09303_),
    .B2(_00192_),
    .Y(_09305_)
  );
  sg13g2_nor2_1 _18911_ (
    .A(_01034_),
    .B(_09305_),
    .Y(_09306_)
  );
  sg13g2_a22oi_1 _18912_ (
    .A1(_09300_),
    .A2(_09301_),
    .B1(_01351_),
    .B2(_09306_),
    .Y(_09307_)
  );
  sg13g2_a21oi_1 _18913_ (
    .A1(_06862_),
    .A2(_02887_),
    .B1(_02990_),
    .Y(_09308_)
  );
  sg13g2_a21oi_1 _18914_ (
    .A1(_06088_),
    .A2(_00878_),
    .B1(addr_i_3_),
    .Y(_09309_)
  );
  sg13g2_or4_1 _18915_ (
    .A(_00268_),
    .B(_05568_),
    .C(_09308_),
    .D(_09309_),
    .X(_09310_)
  );
  sg13g2_nand2_1 _18916_ (
    .A(_02513_),
    .B(_01168_),
    .Y(_09311_)
  );
  sg13g2_a21oi_1 _18917_ (
    .A1(_02694_),
    .A2(_01422_),
    .B1(_00822_),
    .Y(_09312_)
  );
  sg13g2_a21oi_1 _18918_ (
    .A1(_02529_),
    .A2(_03936_),
    .B1(addr_i_5_),
    .Y(_09313_)
  );
  sg13g2_a22oi_1 _18919_ (
    .A1(_01169_),
    .A2(_09311_),
    .B1(_09312_),
    .B2(_09313_),
    .Y(_09314_)
  );
  sg13g2_nor2_1 _18920_ (
    .A(_00290_),
    .B(_09314_),
    .Y(_09316_)
  );
  sg13g2_a21oi_1 _18921_ (
    .A1(_00277_),
    .A2(_09310_),
    .B1(_09316_),
    .Y(_09317_)
  );
  sg13g2_nand2_1 _18922_ (
    .A(addr_i_8_),
    .B(_01024_),
    .Y(_09318_)
  );
  sg13g2_o21ai_1 _18923_ (
    .A1(addr_i_4_),
    .A2(_01928_),
    .B1(_09318_),
    .Y(_09319_)
  );
  sg13g2_nor2_1 _18924_ (
    .A(_06017_),
    .B(_00522_),
    .Y(_09320_)
  );
  sg13g2_a21oi_1 _18925_ (
    .A1(addr_i_3_),
    .A2(_09319_),
    .B1(_09320_),
    .Y(_09321_)
  );
  sg13g2_nor2_1 _18926_ (
    .A(_03886_),
    .B(_01912_),
    .Y(_09322_)
  );
  sg13g2_nand2_1 _18927_ (
    .A(_00711_),
    .B(_00578_),
    .Y(_09323_)
  );
  sg13g2_a21oi_1 _18928_ (
    .A1(_07706_),
    .A2(_09323_),
    .B1(addr_i_5_),
    .Y(_09324_)
  );
  sg13g2_o21ai_1 _18929_ (
    .A1(_09322_),
    .A2(_09324_),
    .B1(_01633_),
    .Y(_09325_)
  );
  sg13g2_o21ai_1 _18930_ (
    .A1(_01543_),
    .A2(_09321_),
    .B1(_09325_),
    .Y(_09327_)
  );
  sg13g2_nor2_1 _18931_ (
    .A(_04661_),
    .B(_04355_),
    .Y(_09328_)
  );
  sg13g2_a21oi_1 _18932_ (
    .A1(_08598_),
    .A2(_02498_),
    .B1(_09328_),
    .Y(_09329_)
  );
  sg13g2_nor3_1 _18933_ (
    .A(_00715_),
    .B(_02424_),
    .C(_00009_),
    .Y(_09330_)
  );
  sg13g2_nor3_1 _18934_ (
    .A(_01920_),
    .B(_01936_),
    .C(_02411_),
    .Y(_09331_)
  );
  sg13g2_nor3_1 _18935_ (
    .A(_00791_),
    .B(_01290_),
    .C(_08951_),
    .Y(_09332_)
  );
  sg13g2_nor4_1 _18936_ (
    .A(addr_i_9_),
    .B(_09330_),
    .C(_09331_),
    .D(_09332_),
    .Y(_09333_)
  );
  sg13g2_o21ai_1 _18937_ (
    .A1(addr_i_3_),
    .A2(_09329_),
    .B1(_09333_),
    .Y(_09334_)
  );
  sg13g2_a21o_1 _18938_ (
    .A1(addr_i_2_),
    .A2(_00412_),
    .B1(_03565_),
    .X(_09335_)
  );
  sg13g2_a21oi_1 _18939_ (
    .A1(_00403_),
    .A2(_00870_),
    .B1(addr_i_4_),
    .Y(_09336_)
  );
  sg13g2_a22oi_1 _18940_ (
    .A1(addr_i_3_),
    .A2(_09335_),
    .B1(_09336_),
    .B2(_00290_),
    .Y(_09338_)
  );
  sg13g2_nor3_1 _18941_ (
    .A(_09327_),
    .B(_09334_),
    .C(_09338_),
    .Y(_09339_)
  );
  sg13g2_a22oi_1 _18942_ (
    .A1(_09307_),
    .A2(_09317_),
    .B1(_09339_),
    .B2(_03841_),
    .Y(_09340_)
  );
  sg13g2_nor2_1 _18943_ (
    .A(addr_i_11_),
    .B(_09340_),
    .Y(_09341_)
  );
  sg13g2_o21ai_1 _18944_ (
    .A1(_00192_),
    .A2(_09094_),
    .B1(addr_i_3_),
    .Y(_09342_)
  );
  sg13g2_a21o_1 _18945_ (
    .A1(_03669_),
    .A2(_06122_),
    .B1(addr_i_2_),
    .X(_09343_)
  );
  sg13g2_nand3_1 _18946_ (
    .A(_01425_),
    .B(_09342_),
    .C(_09343_),
    .Y(_09344_)
  );
  sg13g2_a21oi_1 _18947_ (
    .A1(_02012_),
    .A2(_01007_),
    .B1(addr_i_4_),
    .Y(_09345_)
  );
  sg13g2_a22oi_1 _18948_ (
    .A1(_00910_),
    .A2(_05985_),
    .B1(_09345_),
    .B2(_03577_),
    .Y(_09346_)
  );
  sg13g2_a21oi_1 _18949_ (
    .A1(_03521_),
    .A2(_09346_),
    .B1(_01034_),
    .Y(_09347_)
  );
  sg13g2_nand2_1 _18950_ (
    .A(_01273_),
    .B(_01029_),
    .Y(_09349_)
  );
  sg13g2_a22oi_1 _18951_ (
    .A1(addr_i_5_),
    .A2(_09349_),
    .B1(_03501_),
    .B2(_06276_),
    .Y(_09350_)
  );
  sg13g2_a21oi_1 _18952_ (
    .A1(_04727_),
    .A2(_02965_),
    .B1(_07514_),
    .Y(_09351_)
  );
  sg13g2_o21ai_1 _18953_ (
    .A1(_00060_),
    .A2(_09350_),
    .B1(_09351_),
    .Y(_09352_)
  );
  sg13g2_nand3_1 _18954_ (
    .A(_00322_),
    .B(_01473_),
    .C(_06132_),
    .Y(_09353_)
  );
  sg13g2_nand4_1 _18955_ (
    .A(addr_i_3_),
    .B(_00520_),
    .C(_02479_),
    .D(_00477_),
    .Y(_09354_)
  );
  sg13g2_nand3_1 _18956_ (
    .A(_00276_),
    .B(_09353_),
    .C(_09354_),
    .Y(_09355_)
  );
  sg13g2_nand3_1 _18957_ (
    .A(addr_i_9_),
    .B(_09352_),
    .C(_09355_),
    .Y(_09356_)
  );
  sg13g2_a22oi_1 _18958_ (
    .A1(_01119_),
    .A2(_09344_),
    .B1(_09347_),
    .B2(_09356_),
    .Y(_09357_)
  );
  sg13g2_o21ai_1 _18959_ (
    .A1(_00624_),
    .A2(_00998_),
    .B1(addr_i_4_),
    .Y(_09358_)
  );
  sg13g2_o21ai_1 _18960_ (
    .A1(_09495_),
    .A2(_02321_),
    .B1(addr_i_6_),
    .Y(_09360_)
  );
  sg13g2_and4_1 _18961_ (
    .A(addr_i_2_),
    .B(_08291_),
    .C(_09358_),
    .D(_09360_),
    .X(_09361_)
  );
  sg13g2_a21oi_1 _18962_ (
    .A1(_01786_),
    .A2(_03212_),
    .B1(addr_i_7_),
    .Y(_09362_)
  );
  sg13g2_a22oi_1 _18963_ (
    .A1(addr_i_3_),
    .A2(_00644_),
    .B1(_09362_),
    .B2(addr_i_2_),
    .Y(_09363_)
  );
  sg13g2_o21ai_1 _18964_ (
    .A1(_01519_),
    .A2(_02361_),
    .B1(_06927_),
    .Y(_09364_)
  );
  sg13g2_o21ai_1 _18965_ (
    .A1(_09361_),
    .A2(_09363_),
    .B1(_09364_),
    .Y(_09365_)
  );
  sg13g2_o21ai_1 _18966_ (
    .A1(_08332_),
    .A2(_02462_),
    .B1(addr_i_5_),
    .Y(_09366_)
  );
  sg13g2_a21oi_1 _18967_ (
    .A1(_04384_),
    .A2(_06773_),
    .B1(_05711_),
    .Y(_09367_)
  );
  sg13g2_nor2_1 _18968_ (
    .A(_05237_),
    .B(_09367_),
    .Y(_09368_)
  );
  sg13g2_a22oi_1 _18969_ (
    .A1(_00360_),
    .A2(_09366_),
    .B1(_09368_),
    .B2(addr_i_2_),
    .Y(_09369_)
  );
  sg13g2_o21ai_1 _18970_ (
    .A1(_08056_),
    .A2(_01946_),
    .B1(addr_i_8_),
    .Y(_09372_)
  );
  sg13g2_a21oi_1 _18971_ (
    .A1(_03953_),
    .A2(_00595_),
    .B1(addr_i_4_),
    .Y(_09373_)
  );
  sg13g2_a21oi_1 _18972_ (
    .A1(_09510_),
    .A2(_00789_),
    .B1(_00343_),
    .Y(_09374_)
  );
  sg13g2_a21oi_1 _18973_ (
    .A1(addr_i_3_),
    .A2(_09221_),
    .B1(_01867_),
    .Y(_09375_)
  );
  sg13g2_nor2_1 _18974_ (
    .A(_06154_),
    .B(_09375_),
    .Y(_09376_)
  );
  sg13g2_nor4_1 _18975_ (
    .A(_02344_),
    .B(_09373_),
    .C(_09374_),
    .D(_09376_),
    .Y(_09377_)
  );
  sg13g2_nor3_1 _18976_ (
    .A(_09369_),
    .B(_09372_),
    .C(_09377_),
    .Y(_09378_)
  );
  sg13g2_a22oi_1 _18977_ (
    .A1(_03259_),
    .A2(_09365_),
    .B1(_09378_),
    .B2(addr_i_9_),
    .Y(_09379_)
  );
  sg13g2_or3_1 _18978_ (
    .A(addr_i_10_),
    .B(_09357_),
    .C(_09379_),
    .X(_09380_)
  );
  sg13g2_nor2_1 _18979_ (
    .A(addr_i_3_),
    .B(_01936_),
    .Y(_09381_)
  );
  sg13g2_o21ai_1 _18980_ (
    .A1(addr_i_4_),
    .A2(_06017_),
    .B1(_01928_),
    .Y(_09383_)
  );
  sg13g2_a221oi_1 _18981_ (
    .A1(addr_i_4_),
    .A2(_01537_),
    .B1(addr_i_5_),
    .B2(_09383_),
    .C1(_00535_),
    .Y(_09384_)
  );
  sg13g2_a22oi_1 _18982_ (
    .A1(_05116_),
    .A2(_09381_),
    .B1(_09384_),
    .B2(addr_i_2_),
    .Y(_09385_)
  );
  sg13g2_a22oi_1 _18983_ (
    .A1(addr_i_4_),
    .A2(_03775_),
    .B1(_02542_),
    .B2(_08785_),
    .Y(_09386_)
  );
  sg13g2_a21oi_1 _18984_ (
    .A1(addr_i_2_),
    .A2(_01917_),
    .B1(_00873_),
    .Y(_09387_)
  );
  sg13g2_nor2_1 _18985_ (
    .A(_09386_),
    .B(_09387_),
    .Y(_09388_)
  );
  sg13g2_a22oi_1 _18986_ (
    .A1(_00170_),
    .A2(_00901_),
    .B1(_09385_),
    .B2(_09388_),
    .Y(_09389_)
  );
  sg13g2_o21ai_1 _18987_ (
    .A1(addr_i_6_),
    .A2(_05112_),
    .B1(addr_i_4_),
    .Y(_09390_)
  );
  sg13g2_o21ai_1 _18988_ (
    .A1(_06198_),
    .A2(_05112_),
    .B1(addr_i_6_),
    .Y(_09391_)
  );
  sg13g2_nand2_1 _18989_ (
    .A(_09390_),
    .B(_09391_),
    .Y(_09392_)
  );
  sg13g2_a21oi_1 _18990_ (
    .A1(_05139_),
    .A2(_08349_),
    .B1(addr_i_4_),
    .Y(_09394_)
  );
  sg13g2_a22oi_1 _18991_ (
    .A1(addr_i_8_),
    .A2(_00406_),
    .B1(addr_i_5_),
    .B2(addr_i_6_),
    .Y(_09395_)
  );
  sg13g2_a22oi_1 _18992_ (
    .A1(addr_i_5_),
    .A2(_09392_),
    .B1(_09394_),
    .B2(_09395_),
    .Y(_09396_)
  );
  sg13g2_o21ai_1 _18993_ (
    .A1(_06187_),
    .A2(_05112_),
    .B1(addr_i_5_),
    .Y(_09397_)
  );
  sg13g2_a21oi_1 _18994_ (
    .A1(_08511_),
    .A2(_09397_),
    .B1(addr_i_4_),
    .Y(_09398_)
  );
  sg13g2_a21oi_1 _18995_ (
    .A1(_05902_),
    .A2(_02781_),
    .B1(_01636_),
    .Y(_09399_)
  );
  sg13g2_nor4_1 _18996_ (
    .A(addr_i_3_),
    .B(_01112_),
    .C(_09398_),
    .D(_09399_),
    .Y(_09400_)
  );
  sg13g2_a22oi_1 _18997_ (
    .A1(addr_i_3_),
    .A2(_09396_),
    .B1(_09400_),
    .B2(addr_i_7_),
    .Y(_09401_)
  );
  sg13g2_a21o_1 _18998_ (
    .A1(addr_i_7_),
    .A2(_09389_),
    .B1(_09401_),
    .X(_09402_)
  );
  sg13g2_nand3_1 _18999_ (
    .A(addr_i_3_),
    .B(_00831_),
    .C(_03113_),
    .Y(_09403_)
  );
  sg13g2_a22oi_1 _19000_ (
    .A1(_01420_),
    .A2(_02154_),
    .B1(_09403_),
    .B2(_00377_),
    .Y(_09405_)
  );
  sg13g2_nand2_1 _19001_ (
    .A(_01212_),
    .B(_02406_),
    .Y(_09406_)
  );
  sg13g2_nor3_1 _19002_ (
    .A(addr_i_4_),
    .B(addr_i_7_),
    .C(_05220_),
    .Y(_09407_)
  );
  sg13g2_a22oi_1 _19003_ (
    .A1(addr_i_4_),
    .A2(_09406_),
    .B1(_09407_),
    .B2(addr_i_3_),
    .Y(_09408_)
  );
  sg13g2_a22oi_1 _19004_ (
    .A1(addr_i_7_),
    .A2(_02821_),
    .B1(_00474_),
    .B2(_06695_),
    .Y(_09409_)
  );
  sg13g2_o21ai_1 _19005_ (
    .A1(_09405_),
    .A2(_09408_),
    .B1(_09409_),
    .Y(_09410_)
  );
  sg13g2_o21ai_1 _19006_ (
    .A1(_03523_),
    .A2(_00329_),
    .B1(_00479_),
    .Y(_09411_)
  );
  sg13g2_nand2_1 _19007_ (
    .A(_04650_),
    .B(_09411_),
    .Y(_09412_)
  );
  sg13g2_a22oi_1 _19008_ (
    .A1(_01302_),
    .A2(_04941_),
    .B1(_09412_),
    .B2(_01779_),
    .Y(_09413_)
  );
  sg13g2_a21oi_1 _19009_ (
    .A1(_03022_),
    .A2(_06960_),
    .B1(_03132_),
    .Y(_09414_)
  );
  sg13g2_nor2_1 _19010_ (
    .A(addr_i_6_),
    .B(_00972_),
    .Y(_09416_)
  );
  sg13g2_a21oi_1 _19011_ (
    .A1(addr_i_4_),
    .A2(_02732_),
    .B1(_00697_),
    .Y(_09417_)
  );
  sg13g2_o21ai_1 _19012_ (
    .A1(_00034_),
    .A2(_00482_),
    .B1(_00429_),
    .Y(_09418_)
  );
  sg13g2_a22oi_1 _19013_ (
    .A1(_00771_),
    .A2(_09416_),
    .B1(_09417_),
    .B2(_09418_),
    .Y(_09419_)
  );
  sg13g2_nor4_1 _19014_ (
    .A(addr_i_9_),
    .B(_09413_),
    .C(_09414_),
    .D(_09419_),
    .Y(_09420_)
  );
  sg13g2_a221oi_1 _19015_ (
    .A1(addr_i_9_),
    .A2(_09402_),
    .B1(_09410_),
    .B2(_09420_),
    .C1(addr_i_10_),
    .Y(_09421_)
  );
  sg13g2_a21oi_1 _19016_ (
    .A1(_00914_),
    .A2(_05710_),
    .B1(_06017_),
    .Y(_09422_)
  );
  sg13g2_a21oi_1 _19017_ (
    .A1(_00516_),
    .A2(_03465_),
    .B1(_08464_),
    .Y(_09423_)
  );
  sg13g2_o21ai_1 _19018_ (
    .A1(_09422_),
    .A2(_09423_),
    .B1(_03652_),
    .Y(_09424_)
  );
  sg13g2_nand2_1 _19019_ (
    .A(addr_i_8_),
    .B(_00011_),
    .Y(_09425_)
  );
  sg13g2_o21ai_1 _19020_ (
    .A1(_00284_),
    .A2(_01923_),
    .B1(_09425_),
    .Y(_09427_)
  );
  sg13g2_nand2_1 _19021_ (
    .A(_01019_),
    .B(_09427_),
    .Y(_09428_)
  );
  sg13g2_nand2_1 _19022_ (
    .A(addr_i_3_),
    .B(_05102_),
    .Y(_09429_)
  );
  sg13g2_nand3_1 _19023_ (
    .A(_09424_),
    .B(_09428_),
    .C(_09429_),
    .Y(_09430_)
  );
  sg13g2_a21oi_1 _19024_ (
    .A1(addr_i_3_),
    .A2(_00939_),
    .B1(_01500_),
    .Y(_09431_)
  );
  sg13g2_a21oi_1 _19025_ (
    .A1(_01420_),
    .A2(_03886_),
    .B1(_02008_),
    .Y(_09432_)
  );
  sg13g2_o21ai_1 _19026_ (
    .A1(addr_i_4_),
    .A2(_09431_),
    .B1(_09432_),
    .Y(_09433_)
  );
  sg13g2_o21ai_1 _19027_ (
    .A1(addr_i_4_),
    .A2(_00016_),
    .B1(_01948_),
    .Y(_09434_)
  );
  sg13g2_a21oi_1 _19028_ (
    .A1(_04284_),
    .A2(_02141_),
    .B1(_02152_),
    .Y(_09435_)
  );
  sg13g2_nor2_1 _19029_ (
    .A(_00648_),
    .B(_09435_),
    .Y(_09436_)
  );
  sg13g2_a221oi_1 _19030_ (
    .A1(_02064_),
    .A2(_01998_),
    .B1(_09434_),
    .B2(addr_i_5_),
    .C1(_09436_),
    .Y(_09438_)
  );
  sg13g2_o21ai_1 _19031_ (
    .A1(_01319_),
    .A2(_00110_),
    .B1(addr_i_5_),
    .Y(_09439_)
  );
  sg13g2_o21ai_1 _19032_ (
    .A1(_00165_),
    .A2(_07998_),
    .B1(addr_i_6_),
    .Y(_09440_)
  );
  sg13g2_a21o_1 _19033_ (
    .A1(_09439_),
    .A2(_09440_),
    .B1(addr_i_2_),
    .X(_09441_)
  );
  sg13g2_a21oi_1 _19034_ (
    .A1(_02089_),
    .A2(_01692_),
    .B1(_00145_),
    .Y(_09442_)
  );
  sg13g2_nor2_1 _19035_ (
    .A(_08725_),
    .B(_09442_),
    .Y(_09443_)
  );
  sg13g2_a221oi_1 _19036_ (
    .A1(_02530_),
    .A2(_09438_),
    .B1(_09441_),
    .B2(_09443_),
    .C1(addr_i_8_),
    .Y(_09444_)
  );
  sg13g2_a221oi_1 _19037_ (
    .A1(addr_i_7_),
    .A2(_09430_),
    .B1(_09433_),
    .B2(_01119_),
    .C1(_09444_),
    .Y(_09445_)
  );
  sg13g2_nor2_1 _19038_ (
    .A(_01211_),
    .B(_09445_),
    .Y(_09446_)
  );
  sg13g2_nor3_1 _19039_ (
    .A(_02404_),
    .B(_02322_),
    .C(_02980_),
    .Y(_09447_)
  );
  sg13g2_a22oi_1 _19040_ (
    .A1(_00701_),
    .A2(_00194_),
    .B1(_09447_),
    .B2(addr_i_2_),
    .Y(_09449_)
  );
  sg13g2_a21oi_1 _19041_ (
    .A1(_00069_),
    .A2(_00070_),
    .B1(_01339_),
    .Y(_09450_)
  );
  sg13g2_o21ai_1 _19042_ (
    .A1(_09449_),
    .A2(_09450_),
    .B1(addr_i_6_),
    .Y(_09451_)
  );
  sg13g2_a21oi_1 _19043_ (
    .A1(addr_i_4_),
    .A2(_07570_),
    .B1(_02794_),
    .Y(_09452_)
  );
  sg13g2_nor2_1 _19044_ (
    .A(_09205_),
    .B(_09452_),
    .Y(_09453_)
  );
  sg13g2_a22oi_1 _19045_ (
    .A1(_01194_),
    .A2(_01240_),
    .B1(_09453_),
    .B2(_00367_),
    .Y(_09454_)
  );
  sg13g2_o21ai_1 _19046_ (
    .A1(_02153_),
    .A2(_09506_),
    .B1(_05402_),
    .Y(_09455_)
  );
  sg13g2_a21oi_1 _19047_ (
    .A1(_00220_),
    .A2(_09455_),
    .B1(_00122_),
    .Y(_09456_)
  );
  sg13g2_a22oi_1 _19048_ (
    .A1(_02803_),
    .A2(_01623_),
    .B1(_09456_),
    .B2(addr_i_3_),
    .Y(_09457_)
  );
  sg13g2_nand3_1 _19049_ (
    .A(addr_i_4_),
    .B(addr_i_7_),
    .C(_01656_),
    .Y(_09458_)
  );
  sg13g2_nand3_1 _19050_ (
    .A(addr_i_3_),
    .B(_00353_),
    .C(_09458_),
    .Y(_09460_)
  );
  sg13g2_nand2b_1 _19051_ (
    .A_N(_09457_),
    .B(_09460_),
    .Y(_09461_)
  );
  sg13g2_o21ai_1 _19052_ (
    .A1(_00087_),
    .A2(_02330_),
    .B1(addr_i_4_),
    .Y(_09462_)
  );
  sg13g2_o21ai_1 _19053_ (
    .A1(_07647_),
    .A2(_02639_),
    .B1(addr_i_3_),
    .Y(_09463_)
  );
  sg13g2_nand3_1 _19054_ (
    .A(_01137_),
    .B(_09462_),
    .C(_09463_),
    .Y(_09464_)
  );
  sg13g2_a221oi_1 _19055_ (
    .A1(_01365_),
    .A2(_03572_),
    .B1(_09464_),
    .B2(addr_i_5_),
    .C1(addr_i_8_),
    .Y(_09465_)
  );
  sg13g2_a221oi_1 _19056_ (
    .A1(_09451_),
    .A2(_09454_),
    .B1(_09461_),
    .B2(_09465_),
    .C1(_02221_),
    .Y(_09466_)
  );
  sg13g2_nor4_1 _19057_ (
    .A(_03040_),
    .B(_09421_),
    .C(_09446_),
    .D(_09466_),
    .Y(_09467_)
  );
  sg13g2_a22oi_1 _19058_ (
    .A1(_09341_),
    .A2(_09380_),
    .B1(addr_i_12_),
    .B2(_09467_),
    .Y(_09468_)
  );
  sg13g2_a21o_1 _19059_ (
    .A1(_09283_),
    .A2(_09298_),
    .B1(_09468_),
    .X(data_o_9_)
  );
endmodule
